-- nios2_ht18_lemonde_streit.vhd

-- Generated using ACDS version 13.0sp1 232 at 2018.09.24.13:29:06

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios2_ht18_lemonde_streit is
	port (
		switches18_export  : in    std_logic_vector(17 downto 0) := (others => '0'); --  switches18.export
		keys4_export       : in    std_logic_vector(3 downto 0)  := (others => '0'); --       keys4.export
		leds_red18_export  : out   std_logic_vector(17 downto 0);                    --  leds_red18.export
		leds_green9_export : out   std_logic_vector(8 downto 0);                     -- leds_green9.export
		hex_high28_export  : out   std_logic_vector(27 downto 0);                    --  hex_high28.export
		hex_low28_export   : out   std_logic_vector(27 downto 0);                    --   hex_low28.export
		sdram_wire_addr    : out   std_logic_vector(11 downto 0);                    --  sdram_wire.addr
		sdram_wire_ba      : out   std_logic_vector(1 downto 0);                     --            .ba
		sdram_wire_cas_n   : out   std_logic;                                        --            .cas_n
		sdram_wire_cke     : out   std_logic;                                        --            .cke
		sdram_wire_cs_n    : out   std_logic;                                        --            .cs_n
		sdram_wire_dq      : inout std_logic_vector(15 downto 0) := (others => '0'); --            .dq
		sdram_wire_dqm     : out   std_logic_vector(1 downto 0);                     --            .dqm
		sdram_wire_ras_n   : out   std_logic;                                        --            .ras_n
		sdram_wire_we_n    : out   std_logic;                                        --            .we_n
		clk_clk            : in    std_logic                     := '0';             --         clk.clk
		reset_reset_n      : in    std_logic                     := '0';             --       reset.reset_n
		sdram_clk_clk      : out   std_logic;                                        --   sdram_clk.clk
		sram_wire_DQ       : inout std_logic_vector(15 downto 0) := (others => '0'); --   sram_wire.DQ
		sram_wire_ADDR     : out   std_logic_vector(17 downto 0);                    --            .ADDR
		sram_wire_LB_N     : out   std_logic;                                        --            .LB_N
		sram_wire_UB_N     : out   std_logic;                                        --            .UB_N
		sram_wire_CE_N     : out   std_logic;                                        --            .CE_N
		sram_wire_OE_N     : out   std_logic;                                        --            .OE_N
		sram_wire_WE_N     : out   std_logic                                         --            .WE_N
	);
end entity nios2_ht18_lemonde_streit;

architecture rtl of nios2_ht18_lemonde_streit is
	component nios2_ht18_lemonde_streit_nios2_ht18_lemonde_streit is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(24 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(24 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component nios2_ht18_lemonde_streit_nios2_ht18_lemonde_streit;

	component nios2_ht18_lemonde_streit_onchip_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component nios2_ht18_lemonde_streit_onchip_memory;

	component nios2_ht18_lemonde_streit_ht18_lemonde_streit is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component nios2_ht18_lemonde_streit_ht18_lemonde_streit;

	component nios2_ht18_lemonde_streit_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios2_ht18_lemonde_streit_jtag_uart_0;

	component nios2_ht18_lemonde_streit_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component nios2_ht18_lemonde_streit_timer_0;

	component nios2_ht18_lemonde_streit_timer_1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component nios2_ht18_lemonde_streit_timer_1;

	component nios2_ht18_lemonde_streit_p_counter is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			write         : in  std_logic                     := 'X';             -- write
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component nios2_ht18_lemonde_streit_p_counter;

	component nios2_ht18_lemonde_streit_de2_pio_toggles18 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(17 downto 0) := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component nios2_ht18_lemonde_streit_de2_pio_toggles18;

	component nios2_ht18_lemonde_streit_de2_pio_keys4 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component nios2_ht18_lemonde_streit_de2_pio_keys4;

	component nios2_ht18_lemonde_streit_de2_pio_redled18 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(17 downto 0)                     -- export
		);
	end component nios2_ht18_lemonde_streit_de2_pio_redled18;

	component nios2_ht18_lemonde_streit_de2_pio_greenled9 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(8 downto 0)                      -- export
		);
	end component nios2_ht18_lemonde_streit_de2_pio_greenled9;

	component nios2_ht18_lemonde_streit_de2_pio_hex_high28 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(27 downto 0)                     -- export
		);
	end component nios2_ht18_lemonde_streit_de2_pio_hex_high28;

	component nios2_ht18_lemonde_streit_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component nios2_ht18_lemonde_streit_sdram;

	component nios2_ht18_lemonde_streit_up_clocks_0 is
		port (
			CLOCK_50    : in  std_logic := 'X'; -- clk
			reset       : in  std_logic := 'X'; -- reset
			sys_clk     : out std_logic;        -- clk
			sys_reset_n : out std_logic;        -- reset_n
			SDRAM_CLK   : out std_logic         -- clk
		);
	end component nios2_ht18_lemonde_streit_up_clocks_0;

	component nios2_ht18_lemonde_streit_sram is
		port (
			clk           : in    std_logic                     := 'X';             -- clk
			reset         : in    std_logic                     := 'X';             -- reset
			SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			SRAM_ADDR     : out   std_logic_vector(17 downto 0);                    -- export
			SRAM_LB_N     : out   std_logic;                                        -- export
			SRAM_UB_N     : out   std_logic;                                        -- export
			SRAM_CE_N     : out   std_logic;                                        -- export
			SRAM_OE_N     : out   std_logic;                                        -- export
			SRAM_WE_N     : out   std_logic;                                        -- export
			address       : in    std_logic_vector(17 downto 0) := (others => 'X'); -- address
			byteenable    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			read          : in    std_logic                     := 'X';             -- read
			write         : in    std_logic                     := 'X';             -- write
			writedata     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out   std_logic_vector(15 downto 0);                    -- readdata
			readdatavalid : out   std_logic                                         -- readdatavalid
		);
	end component nios2_ht18_lemonde_streit_sram;

	component altera_merlin_master_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(99 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component altera_merlin_master_agent;

	component nios2_ht18_lemonde_streit_addr_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(99 downto 0);                    -- data
			src_channel        : out std_logic_vector(14 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios2_ht18_lemonde_streit_addr_router;

	component nios2_ht18_lemonde_streit_addr_router_001 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(99 downto 0);                    -- data
			src_channel        : out std_logic_vector(14 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios2_ht18_lemonde_streit_addr_router_001;

	component nios2_ht18_lemonde_streit_id_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(99 downto 0);                    -- data
			src_channel        : out std_logic_vector(14 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios2_ht18_lemonde_streit_id_router;

	component nios2_ht18_lemonde_streit_id_router_001 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(99 downto 0);                    -- data
			src_channel        : out std_logic_vector(14 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios2_ht18_lemonde_streit_id_router_001;

	component nios2_ht18_lemonde_streit_id_router_013 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(81 downto 0);                    -- data
			src_channel        : out std_logic_vector(14 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios2_ht18_lemonde_streit_id_router_013;

	component altera_merlin_burst_adapter is
		generic (
			PKT_ADDR_H                : integer := 79;
			PKT_ADDR_L                : integer := 48;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BYTE_CNT_H            : integer := 5;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 83;
			PKT_BYTEEN_L              : integer := 80;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 88;
			PKT_BURST_TYPE_L          : integer := 87;
			PKT_BURSTWRAP_H           : integer := 11;
			PKT_BURSTWRAP_L           : integer := 6;
			PKT_TRANS_COMPRESSED_READ : integer := 14;
			PKT_TRANS_WRITE           : integer := 13;
			PKT_TRANS_READ            : integer := 12;
			OUT_NARROW_SIZE           : integer := 0;
			IN_NARROW_SIZE            : integer := 0;
			OUT_FIXED                 : integer := 0;
			OUT_COMPLETE_WRAP         : integer := 0;
			ST_DATA_W                 : integer := 89;
			ST_CHANNEL_W              : integer := 8;
			OUT_BYTE_CNT_H            : integer := 5;
			OUT_BURSTWRAP_H           : integer := 11;
			COMPRESSED_READ_SUPPORT   : integer := 1;
			BYTEENABLE_SYNTHESIS      : integer := 0;
			PIPE_INPUTS               : integer := 0;
			NO_WRAP_SUPPORT           : integer := 0;
			BURSTWRAP_CONST_MASK      : integer := 0;
			BURSTWRAP_CONST_VALUE     : integer := -1
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			sink0_valid           : in  std_logic                     := 'X';             -- valid
			sink0_data            : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                        -- ready
			source0_valid         : out std_logic;                                        -- valid
			source0_data          : out std_logic_vector(81 downto 0);                    -- data
			source0_channel       : out std_logic_vector(14 downto 0);                    -- channel
			source0_startofpacket : out std_logic;                                        -- startofpacket
			source0_endofpacket   : out std_logic;                                        -- endofpacket
			source0_ready         : in  std_logic                     := 'X'              -- ready
		);
	end component altera_merlin_burst_adapter;

	component nios2_ht18_lemonde_streit_cmd_xbar_demux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			sink_ready          : out std_logic;                                        -- ready
			sink_channel        : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink_valid          : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready          : in  std_logic                     := 'X';             -- ready
			src0_valid          : out std_logic;                                        -- valid
			src0_data           : out std_logic_vector(99 downto 0);                    -- data
			src0_channel        : out std_logic_vector(14 downto 0);                    -- channel
			src0_startofpacket  : out std_logic;                                        -- startofpacket
			src0_endofpacket    : out std_logic;                                        -- endofpacket
			src1_ready          : in  std_logic                     := 'X';             -- ready
			src1_valid          : out std_logic;                                        -- valid
			src1_data           : out std_logic_vector(99 downto 0);                    -- data
			src1_channel        : out std_logic_vector(14 downto 0);                    -- channel
			src1_startofpacket  : out std_logic;                                        -- startofpacket
			src1_endofpacket    : out std_logic;                                        -- endofpacket
			src2_ready          : in  std_logic                     := 'X';             -- ready
			src2_valid          : out std_logic;                                        -- valid
			src2_data           : out std_logic_vector(99 downto 0);                    -- data
			src2_channel        : out std_logic_vector(14 downto 0);                    -- channel
			src2_startofpacket  : out std_logic;                                        -- startofpacket
			src2_endofpacket    : out std_logic;                                        -- endofpacket
			src3_ready          : in  std_logic                     := 'X';             -- ready
			src3_valid          : out std_logic;                                        -- valid
			src3_data           : out std_logic_vector(99 downto 0);                    -- data
			src3_channel        : out std_logic_vector(14 downto 0);                    -- channel
			src3_startofpacket  : out std_logic;                                        -- startofpacket
			src3_endofpacket    : out std_logic;                                        -- endofpacket
			src4_ready          : in  std_logic                     := 'X';             -- ready
			src4_valid          : out std_logic;                                        -- valid
			src4_data           : out std_logic_vector(99 downto 0);                    -- data
			src4_channel        : out std_logic_vector(14 downto 0);                    -- channel
			src4_startofpacket  : out std_logic;                                        -- startofpacket
			src4_endofpacket    : out std_logic;                                        -- endofpacket
			src5_ready          : in  std_logic                     := 'X';             -- ready
			src5_valid          : out std_logic;                                        -- valid
			src5_data           : out std_logic_vector(99 downto 0);                    -- data
			src5_channel        : out std_logic_vector(14 downto 0);                    -- channel
			src5_startofpacket  : out std_logic;                                        -- startofpacket
			src5_endofpacket    : out std_logic;                                        -- endofpacket
			src6_ready          : in  std_logic                     := 'X';             -- ready
			src6_valid          : out std_logic;                                        -- valid
			src6_data           : out std_logic_vector(99 downto 0);                    -- data
			src6_channel        : out std_logic_vector(14 downto 0);                    -- channel
			src6_startofpacket  : out std_logic;                                        -- startofpacket
			src6_endofpacket    : out std_logic;                                        -- endofpacket
			src7_ready          : in  std_logic                     := 'X';             -- ready
			src7_valid          : out std_logic;                                        -- valid
			src7_data           : out std_logic_vector(99 downto 0);                    -- data
			src7_channel        : out std_logic_vector(14 downto 0);                    -- channel
			src7_startofpacket  : out std_logic;                                        -- startofpacket
			src7_endofpacket    : out std_logic;                                        -- endofpacket
			src8_ready          : in  std_logic                     := 'X';             -- ready
			src8_valid          : out std_logic;                                        -- valid
			src8_data           : out std_logic_vector(99 downto 0);                    -- data
			src8_channel        : out std_logic_vector(14 downto 0);                    -- channel
			src8_startofpacket  : out std_logic;                                        -- startofpacket
			src8_endofpacket    : out std_logic;                                        -- endofpacket
			src9_ready          : in  std_logic                     := 'X';             -- ready
			src9_valid          : out std_logic;                                        -- valid
			src9_data           : out std_logic_vector(99 downto 0);                    -- data
			src9_channel        : out std_logic_vector(14 downto 0);                    -- channel
			src9_startofpacket  : out std_logic;                                        -- startofpacket
			src9_endofpacket    : out std_logic;                                        -- endofpacket
			src10_ready         : in  std_logic                     := 'X';             -- ready
			src10_valid         : out std_logic;                                        -- valid
			src10_data          : out std_logic_vector(99 downto 0);                    -- data
			src10_channel       : out std_logic_vector(14 downto 0);                    -- channel
			src10_startofpacket : out std_logic;                                        -- startofpacket
			src10_endofpacket   : out std_logic;                                        -- endofpacket
			src11_ready         : in  std_logic                     := 'X';             -- ready
			src11_valid         : out std_logic;                                        -- valid
			src11_data          : out std_logic_vector(99 downto 0);                    -- data
			src11_channel       : out std_logic_vector(14 downto 0);                    -- channel
			src11_startofpacket : out std_logic;                                        -- startofpacket
			src11_endofpacket   : out std_logic;                                        -- endofpacket
			src12_ready         : in  std_logic                     := 'X';             -- ready
			src12_valid         : out std_logic;                                        -- valid
			src12_data          : out std_logic_vector(99 downto 0);                    -- data
			src12_channel       : out std_logic_vector(14 downto 0);                    -- channel
			src12_startofpacket : out std_logic;                                        -- startofpacket
			src12_endofpacket   : out std_logic;                                        -- endofpacket
			src13_ready         : in  std_logic                     := 'X';             -- ready
			src13_valid         : out std_logic;                                        -- valid
			src13_data          : out std_logic_vector(99 downto 0);                    -- data
			src13_channel       : out std_logic_vector(14 downto 0);                    -- channel
			src13_startofpacket : out std_logic;                                        -- startofpacket
			src13_endofpacket   : out std_logic;                                        -- endofpacket
			src14_ready         : in  std_logic                     := 'X';             -- ready
			src14_valid         : out std_logic;                                        -- valid
			src14_data          : out std_logic_vector(99 downto 0);                    -- data
			src14_channel       : out std_logic_vector(14 downto 0);                    -- channel
			src14_startofpacket : out std_logic;                                        -- startofpacket
			src14_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component nios2_ht18_lemonde_streit_cmd_xbar_demux;

	component nios2_ht18_lemonde_streit_cmd_xbar_demux_001 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(99 downto 0);                    -- data
			src0_channel       : out std_logic_vector(14 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(99 downto 0);                    -- data
			src1_channel       : out std_logic_vector(14 downto 0);                    -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic;                                        -- endofpacket
			src2_ready         : in  std_logic                     := 'X';             -- ready
			src2_valid         : out std_logic;                                        -- valid
			src2_data          : out std_logic_vector(99 downto 0);                    -- data
			src2_channel       : out std_logic_vector(14 downto 0);                    -- channel
			src2_startofpacket : out std_logic;                                        -- startofpacket
			src2_endofpacket   : out std_logic;                                        -- endofpacket
			src3_ready         : in  std_logic                     := 'X';             -- ready
			src3_valid         : out std_logic;                                        -- valid
			src3_data          : out std_logic_vector(99 downto 0);                    -- data
			src3_channel       : out std_logic_vector(14 downto 0);                    -- channel
			src3_startofpacket : out std_logic;                                        -- startofpacket
			src3_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component nios2_ht18_lemonde_streit_cmd_xbar_demux_001;

	component nios2_ht18_lemonde_streit_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(99 downto 0);                    -- data
			src_channel         : out std_logic_vector(14 downto 0);                    -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component nios2_ht18_lemonde_streit_cmd_xbar_mux;

	component nios2_ht18_lemonde_streit_rsp_xbar_demux is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(99 downto 0);                    -- data
			src0_channel       : out std_logic_vector(14 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(99 downto 0);                    -- data
			src1_channel       : out std_logic_vector(14 downto 0);                    -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component nios2_ht18_lemonde_streit_rsp_xbar_demux;

	component nios2_ht18_lemonde_streit_rsp_xbar_demux_001 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(99 downto 0);                    -- data
			src0_channel       : out std_logic_vector(14 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component nios2_ht18_lemonde_streit_rsp_xbar_demux_001;

	component nios2_ht18_lemonde_streit_rsp_xbar_mux is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			src_ready            : in  std_logic                     := 'X';             -- ready
			src_valid            : out std_logic;                                        -- valid
			src_data             : out std_logic_vector(99 downto 0);                    -- data
			src_channel          : out std_logic_vector(14 downto 0);                    -- channel
			src_startofpacket    : out std_logic;                                        -- startofpacket
			src_endofpacket      : out std_logic;                                        -- endofpacket
			sink0_ready          : out std_logic;                                        -- ready
			sink0_valid          : in  std_logic                     := 'X';             -- valid
			sink0_channel        : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink0_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready          : out std_logic;                                        -- ready
			sink1_valid          : in  std_logic                     := 'X';             -- valid
			sink1_channel        : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink1_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink1_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready          : out std_logic;                                        -- ready
			sink2_valid          : in  std_logic                     := 'X';             -- valid
			sink2_channel        : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink2_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink2_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready          : out std_logic;                                        -- ready
			sink3_valid          : in  std_logic                     := 'X';             -- valid
			sink3_channel        : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink3_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink3_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink4_ready          : out std_logic;                                        -- ready
			sink4_valid          : in  std_logic                     := 'X';             -- valid
			sink4_channel        : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink4_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink4_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink4_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink5_ready          : out std_logic;                                        -- ready
			sink5_valid          : in  std_logic                     := 'X';             -- valid
			sink5_channel        : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink5_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink5_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink5_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink6_ready          : out std_logic;                                        -- ready
			sink6_valid          : in  std_logic                     := 'X';             -- valid
			sink6_channel        : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink6_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink6_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink6_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink7_ready          : out std_logic;                                        -- ready
			sink7_valid          : in  std_logic                     := 'X';             -- valid
			sink7_channel        : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink7_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink7_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink7_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink8_ready          : out std_logic;                                        -- ready
			sink8_valid          : in  std_logic                     := 'X';             -- valid
			sink8_channel        : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink8_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink8_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink8_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink9_ready          : out std_logic;                                        -- ready
			sink9_valid          : in  std_logic                     := 'X';             -- valid
			sink9_channel        : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink9_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink9_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink9_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink10_ready         : out std_logic;                                        -- ready
			sink10_valid         : in  std_logic                     := 'X';             -- valid
			sink10_channel       : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink10_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink10_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink10_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink11_ready         : out std_logic;                                        -- ready
			sink11_valid         : in  std_logic                     := 'X';             -- valid
			sink11_channel       : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink11_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink11_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink11_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink12_ready         : out std_logic;                                        -- ready
			sink12_valid         : in  std_logic                     := 'X';             -- valid
			sink12_channel       : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink12_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink12_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink12_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink13_ready         : out std_logic;                                        -- ready
			sink13_valid         : in  std_logic                     := 'X';             -- valid
			sink13_channel       : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink13_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink13_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink13_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink14_ready         : out std_logic;                                        -- ready
			sink14_valid         : in  std_logic                     := 'X';             -- valid
			sink14_channel       : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink14_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink14_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink14_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component nios2_ht18_lemonde_streit_rsp_xbar_mux;

	component nios2_ht18_lemonde_streit_rsp_xbar_mux_001 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(99 downto 0);                    -- data
			src_channel         : out std_logic_vector(14 downto 0);                    -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                        -- ready
			sink2_valid         : in  std_logic                     := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready         : out std_logic;                                        -- ready
			sink3_valid         : in  std_logic                     := 'X';             -- valid
			sink3_channel       : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			sink3_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink3_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component nios2_ht18_lemonde_streit_rsp_xbar_mux_001;

	component nios2_ht18_lemonde_streit_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios2_ht18_lemonde_streit_irq_mapper;

	component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(100 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic;                                         -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- address
			csr_read          : in  std_logic                      := 'X';             -- read
			csr_write         : in  std_logic                      := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                     -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                         -- data
			almost_empty_data : out std_logic;                                         -- data
			in_empty          : in  std_logic                      := 'X';             -- empty
			out_empty         : out std_logic;                                         -- empty
			in_error          : in  std_logic                      := 'X';             -- error
			out_error         : out std_logic;                                         -- error
			in_channel        : in  std_logic                      := 'X';             -- channel
			out_channel       : out std_logic                                          -- channel
		);
	end component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component nios2_ht18_lemonde_streit_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(82 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(82 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component nios2_ht18_lemonde_streit_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component nios2_ht18_lemonde_streit_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			out_data          : out std_logic_vector(17 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component nios2_ht18_lemonde_streit_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(99 downto 0);                     -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(99 downto 0)  := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(14 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(100 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                         -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                      := 'X'              -- writeresponsevalid
		);
	end component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent;

	component nios2_ht18_lemonde_streit_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(1 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(81 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(82 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(82 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(17 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2_ht18_lemonde_streit_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent;

	component nios2_ht18_lemonde_streit_width_adapter is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			in_valid             : in  std_logic                     := 'X';             -- valid
			in_channel           : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                     := 'X';             -- endofpacket
			in_ready             : out std_logic;                                        -- ready
			in_data              : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                        -- endofpacket
			out_data             : out std_logic_vector(81 downto 0);                    -- data
			out_channel          : out std_logic_vector(14 downto 0);                    -- channel
			out_valid            : out std_logic;                                        -- valid
			out_ready            : in  std_logic                     := 'X';             -- ready
			out_startofpacket    : out std_logic;                                        -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- data
		);
	end component nios2_ht18_lemonde_streit_width_adapter;

	component nios2_ht18_lemonde_streit_width_adapter_001 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			in_valid             : in  std_logic                     := 'X';             -- valid
			in_channel           : in  std_logic_vector(14 downto 0) := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                     := 'X';             -- endofpacket
			in_ready             : out std_logic;                                        -- ready
			in_data              : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                        -- endofpacket
			out_data             : out std_logic_vector(99 downto 0);                    -- data
			out_channel          : out std_logic_vector(14 downto 0);                    -- channel
			out_valid            : out std_logic;                                        -- valid
			out_ready            : in  std_logic                     := 'X';             -- ready
			out_startofpacket    : out std_logic;                                        -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- data
		);
	end component nios2_ht18_lemonde_streit_width_adapter_001;

	component nios2_ht18_lemonde_streit_nios2_ht18_lemonde_streit_data_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(24 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component nios2_ht18_lemonde_streit_nios2_ht18_lemonde_streit_data_master_translator;

	component nios2_ht18_lemonde_streit_nios2_ht18_lemonde_streit_instruction_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(24 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component nios2_ht18_lemonde_streit_nios2_ht18_lemonde_streit_instruction_master_translator;

	component nios2_ht18_lemonde_streit_onchip_memory_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(12 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2_ht18_lemonde_streit_onchip_memory_s1_translator;

	component nios2_ht18_lemonde_streit_ht18_lemonde_streit_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2_ht18_lemonde_streit_ht18_lemonde_streit_control_slave_translator;

	component nios2_ht18_lemonde_streit_jtag_uart_0_avalon_jtag_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2_ht18_lemonde_streit_jtag_uart_0_avalon_jtag_slave_translator;

	component nios2_ht18_lemonde_streit_nios2_ht18_lemonde_streit_jtag_debug_module_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(8 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2_ht18_lemonde_streit_nios2_ht18_lemonde_streit_jtag_debug_module_translator;

	component nios2_ht18_lemonde_streit_timer_0_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(2 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2_ht18_lemonde_streit_timer_0_s1_translator;

	component nios2_ht18_lemonde_streit_p_counter_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(4 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_read                  : out std_logic;                                        -- read
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2_ht18_lemonde_streit_p_counter_control_slave_translator;

	component nios2_ht18_lemonde_streit_de2_pio_toggles18_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2_ht18_lemonde_streit_de2_pio_toggles18_s1_translator;

	component nios2_ht18_lemonde_streit_sram_avalon_sram_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(17 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(1 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(1 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2_ht18_lemonde_streit_sram_avalon_sram_slave_translator;

	component nios2_ht18_lemonde_streit_sdram_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(21 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(1 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_writebyteenable       : out std_logic_vector(1 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2_ht18_lemonde_streit_sdram_s1_translator;

	component nios2_ht18_lemonde_streit_rst_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			reset_in1  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component nios2_ht18_lemonde_streit_rst_controller;

	component nios2_ht18_lemonde_streit_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component nios2_ht18_lemonde_streit_rst_controller_001;

	component nios2_ht18_lemonde_streit_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			reset_in1  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component nios2_ht18_lemonde_streit_rst_controller_002;

	signal up_clocks_0_sys_clk_clk                                                                                          : std_logic;                      -- up_clocks_0:sys_clk -> [addr_router:clk, addr_router_001:clk, burst_adapter:clk, burst_adapter_001:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_mux:clk, cmd_xbar_mux_003:clk, cmd_xbar_mux_013:clk, cmd_xbar_mux_014:clk, de2_pio_greenled9:clk, de2_pio_greenled9_s1_translator:clk, de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:clk, de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, de2_pio_hex_high28:clk, de2_pio_hex_high28_s1_translator:clk, de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:clk, de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, de2_pio_hex_low28:clk, de2_pio_hex_low28_s1_translator:clk, de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:clk, de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, de2_pio_keys4:clk, de2_pio_keys4_s1_translator:clk, de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:clk, de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, de2_pio_redled18:clk, de2_pio_redled18_s1_translator:clk, de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:clk, de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, de2_pio_toggles18:clk, de2_pio_toggles18_s1_translator:clk, de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:clk, de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, ht18_lemonde_streit:clock, ht18_lemonde_streit_control_slave_translator:clk, ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:clk, ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, irq_mapper:clk, jtag_uart_0:clk, jtag_uart_0_avalon_jtag_slave_translator:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, nios2_ht18_lemonde_streit:clk, nios2_ht18_lemonde_streit_data_master_translator:clk, nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:clk, nios2_ht18_lemonde_streit_instruction_master_translator:clk, nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_ht18_lemonde_streit_jtag_debug_module_translator:clk, nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, onchip_memory:clk, onchip_memory_s1_translator:clk, onchip_memory_s1_translator_avalon_universal_slave_0_agent:clk, onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, p_counter:clk, p_counter_control_slave_translator:clk, p_counter_control_slave_translator_avalon_universal_slave_0_agent:clk, p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller:clk, rst_controller_001:clk, sdram:clk, sdram_s1_translator:clk, sdram_s1_translator_avalon_universal_slave_0_agent:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sram:clk, sram_avalon_sram_slave_translator:clk, sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:clk, sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer_0:clk, timer_0_s1_translator:clk, timer_0_s1_translator_avalon_universal_slave_0_agent:clk, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer_1:clk, timer_1_s1_translator:clk, timer_1_s1_translator_avalon_universal_slave_0_agent:clk, timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk]
	signal nios2_ht18_lemonde_streit_data_master_waitrequest                                                                : std_logic;                      -- nios2_ht18_lemonde_streit_data_master_translator:av_waitrequest -> nios2_ht18_lemonde_streit:d_waitrequest
	signal nios2_ht18_lemonde_streit_data_master_writedata                                                                  : std_logic_vector(31 downto 0);  -- nios2_ht18_lemonde_streit:d_writedata -> nios2_ht18_lemonde_streit_data_master_translator:av_writedata
	signal nios2_ht18_lemonde_streit_data_master_address                                                                    : std_logic_vector(24 downto 0);  -- nios2_ht18_lemonde_streit:d_address -> nios2_ht18_lemonde_streit_data_master_translator:av_address
	signal nios2_ht18_lemonde_streit_data_master_write                                                                      : std_logic;                      -- nios2_ht18_lemonde_streit:d_write -> nios2_ht18_lemonde_streit_data_master_translator:av_write
	signal nios2_ht18_lemonde_streit_data_master_read                                                                       : std_logic;                      -- nios2_ht18_lemonde_streit:d_read -> nios2_ht18_lemonde_streit_data_master_translator:av_read
	signal nios2_ht18_lemonde_streit_data_master_readdata                                                                   : std_logic_vector(31 downto 0);  -- nios2_ht18_lemonde_streit_data_master_translator:av_readdata -> nios2_ht18_lemonde_streit:d_readdata
	signal nios2_ht18_lemonde_streit_data_master_debugaccess                                                                : std_logic;                      -- nios2_ht18_lemonde_streit:jtag_debug_module_debugaccess_to_roms -> nios2_ht18_lemonde_streit_data_master_translator:av_debugaccess
	signal nios2_ht18_lemonde_streit_data_master_byteenable                                                                 : std_logic_vector(3 downto 0);   -- nios2_ht18_lemonde_streit:d_byteenable -> nios2_ht18_lemonde_streit_data_master_translator:av_byteenable
	signal nios2_ht18_lemonde_streit_instruction_master_waitrequest                                                         : std_logic;                      -- nios2_ht18_lemonde_streit_instruction_master_translator:av_waitrequest -> nios2_ht18_lemonde_streit:i_waitrequest
	signal nios2_ht18_lemonde_streit_instruction_master_address                                                             : std_logic_vector(24 downto 0);  -- nios2_ht18_lemonde_streit:i_address -> nios2_ht18_lemonde_streit_instruction_master_translator:av_address
	signal nios2_ht18_lemonde_streit_instruction_master_read                                                                : std_logic;                      -- nios2_ht18_lemonde_streit:i_read -> nios2_ht18_lemonde_streit_instruction_master_translator:av_read
	signal nios2_ht18_lemonde_streit_instruction_master_readdata                                                            : std_logic_vector(31 downto 0);  -- nios2_ht18_lemonde_streit_instruction_master_translator:av_readdata -> nios2_ht18_lemonde_streit:i_readdata
	signal onchip_memory_s1_translator_avalon_anti_slave_0_writedata                                                        : std_logic_vector(31 downto 0);  -- onchip_memory_s1_translator:av_writedata -> onchip_memory:writedata
	signal onchip_memory_s1_translator_avalon_anti_slave_0_address                                                          : std_logic_vector(12 downto 0);  -- onchip_memory_s1_translator:av_address -> onchip_memory:address
	signal onchip_memory_s1_translator_avalon_anti_slave_0_chipselect                                                       : std_logic;                      -- onchip_memory_s1_translator:av_chipselect -> onchip_memory:chipselect
	signal onchip_memory_s1_translator_avalon_anti_slave_0_clken                                                            : std_logic;                      -- onchip_memory_s1_translator:av_clken -> onchip_memory:clken
	signal onchip_memory_s1_translator_avalon_anti_slave_0_write                                                            : std_logic;                      -- onchip_memory_s1_translator:av_write -> onchip_memory:write
	signal onchip_memory_s1_translator_avalon_anti_slave_0_readdata                                                         : std_logic_vector(31 downto 0);  -- onchip_memory:readdata -> onchip_memory_s1_translator:av_readdata
	signal onchip_memory_s1_translator_avalon_anti_slave_0_byteenable                                                       : std_logic_vector(3 downto 0);   -- onchip_memory_s1_translator:av_byteenable -> onchip_memory:byteenable
	signal ht18_lemonde_streit_control_slave_translator_avalon_anti_slave_0_address                                         : std_logic_vector(0 downto 0);   -- ht18_lemonde_streit_control_slave_translator:av_address -> ht18_lemonde_streit:address
	signal ht18_lemonde_streit_control_slave_translator_avalon_anti_slave_0_readdata                                        : std_logic_vector(31 downto 0);  -- ht18_lemonde_streit:readdata -> ht18_lemonde_streit_control_slave_translator:av_readdata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest                                         : std_logic;                      -- jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata                                           : std_logic_vector(31 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address                                             : std_logic_vector(0 downto 0);   -- jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                                          : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write                                               : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write:in
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read                                                : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read:in
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata                                            : std_logic_vector(31 downto 0);  -- jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest                           : std_logic;                      -- nios2_ht18_lemonde_streit:jtag_debug_module_waitrequest -> nios2_ht18_lemonde_streit_jtag_debug_module_translator:av_waitrequest
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0);  -- nios2_ht18_lemonde_streit_jtag_debug_module_translator:av_writedata -> nios2_ht18_lemonde_streit:jtag_debug_module_writedata
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_address                               : std_logic_vector(8 downto 0);   -- nios2_ht18_lemonde_streit_jtag_debug_module_translator:av_address -> nios2_ht18_lemonde_streit:jtag_debug_module_address
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_write                                 : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator:av_write -> nios2_ht18_lemonde_streit:jtag_debug_module_write
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_read                                  : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator:av_read -> nios2_ht18_lemonde_streit:jtag_debug_module_read
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0);  -- nios2_ht18_lemonde_streit:jtag_debug_module_readdata -> nios2_ht18_lemonde_streit_jtag_debug_module_translator:av_readdata
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                           : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator:av_debugaccess -> nios2_ht18_lemonde_streit:jtag_debug_module_debugaccess
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_byteenable                            : std_logic_vector(3 downto 0);   -- nios2_ht18_lemonde_streit_jtag_debug_module_translator:av_byteenable -> nios2_ht18_lemonde_streit:jtag_debug_module_byteenable
	signal timer_0_s1_translator_avalon_anti_slave_0_writedata                                                              : std_logic_vector(15 downto 0);  -- timer_0_s1_translator:av_writedata -> timer_0:writedata
	signal timer_0_s1_translator_avalon_anti_slave_0_address                                                                : std_logic_vector(2 downto 0);   -- timer_0_s1_translator:av_address -> timer_0:address
	signal timer_0_s1_translator_avalon_anti_slave_0_chipselect                                                             : std_logic;                      -- timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	signal timer_0_s1_translator_avalon_anti_slave_0_write                                                                  : std_logic;                      -- timer_0_s1_translator:av_write -> timer_0_s1_translator_avalon_anti_slave_0_write:in
	signal timer_0_s1_translator_avalon_anti_slave_0_readdata                                                               : std_logic_vector(15 downto 0);  -- timer_0:readdata -> timer_0_s1_translator:av_readdata
	signal timer_1_s1_translator_avalon_anti_slave_0_writedata                                                              : std_logic_vector(15 downto 0);  -- timer_1_s1_translator:av_writedata -> timer_1:writedata
	signal timer_1_s1_translator_avalon_anti_slave_0_address                                                                : std_logic_vector(2 downto 0);   -- timer_1_s1_translator:av_address -> timer_1:address
	signal timer_1_s1_translator_avalon_anti_slave_0_chipselect                                                             : std_logic;                      -- timer_1_s1_translator:av_chipselect -> timer_1:chipselect
	signal timer_1_s1_translator_avalon_anti_slave_0_write                                                                  : std_logic;                      -- timer_1_s1_translator:av_write -> timer_1_s1_translator_avalon_anti_slave_0_write:in
	signal timer_1_s1_translator_avalon_anti_slave_0_readdata                                                               : std_logic_vector(15 downto 0);  -- timer_1:readdata -> timer_1_s1_translator:av_readdata
	signal p_counter_control_slave_translator_avalon_anti_slave_0_writedata                                                 : std_logic_vector(31 downto 0);  -- p_counter_control_slave_translator:av_writedata -> p_counter:writedata
	signal p_counter_control_slave_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(4 downto 0);   -- p_counter_control_slave_translator:av_address -> p_counter:address
	signal p_counter_control_slave_translator_avalon_anti_slave_0_write                                                     : std_logic;                      -- p_counter_control_slave_translator:av_write -> p_counter:write
	signal p_counter_control_slave_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(31 downto 0);  -- p_counter:readdata -> p_counter_control_slave_translator:av_readdata
	signal p_counter_control_slave_translator_avalon_anti_slave_0_begintransfer                                             : std_logic;                      -- p_counter_control_slave_translator:av_begintransfer -> p_counter:begintransfer
	signal de2_pio_toggles18_s1_translator_avalon_anti_slave_0_writedata                                                    : std_logic_vector(31 downto 0);  -- de2_pio_toggles18_s1_translator:av_writedata -> de2_pio_toggles18:writedata
	signal de2_pio_toggles18_s1_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(1 downto 0);   -- de2_pio_toggles18_s1_translator:av_address -> de2_pio_toggles18:address
	signal de2_pio_toggles18_s1_translator_avalon_anti_slave_0_chipselect                                                   : std_logic;                      -- de2_pio_toggles18_s1_translator:av_chipselect -> de2_pio_toggles18:chipselect
	signal de2_pio_toggles18_s1_translator_avalon_anti_slave_0_write                                                        : std_logic;                      -- de2_pio_toggles18_s1_translator:av_write -> de2_pio_toggles18_s1_translator_avalon_anti_slave_0_write:in
	signal de2_pio_toggles18_s1_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(31 downto 0);  -- de2_pio_toggles18:readdata -> de2_pio_toggles18_s1_translator:av_readdata
	signal de2_pio_keys4_s1_translator_avalon_anti_slave_0_writedata                                                        : std_logic_vector(31 downto 0);  -- de2_pio_keys4_s1_translator:av_writedata -> de2_pio_keys4:writedata
	signal de2_pio_keys4_s1_translator_avalon_anti_slave_0_address                                                          : std_logic_vector(1 downto 0);   -- de2_pio_keys4_s1_translator:av_address -> de2_pio_keys4:address
	signal de2_pio_keys4_s1_translator_avalon_anti_slave_0_chipselect                                                       : std_logic;                      -- de2_pio_keys4_s1_translator:av_chipselect -> de2_pio_keys4:chipselect
	signal de2_pio_keys4_s1_translator_avalon_anti_slave_0_write                                                            : std_logic;                      -- de2_pio_keys4_s1_translator:av_write -> de2_pio_keys4_s1_translator_avalon_anti_slave_0_write:in
	signal de2_pio_keys4_s1_translator_avalon_anti_slave_0_readdata                                                         : std_logic_vector(31 downto 0);  -- de2_pio_keys4:readdata -> de2_pio_keys4_s1_translator:av_readdata
	signal de2_pio_redled18_s1_translator_avalon_anti_slave_0_writedata                                                     : std_logic_vector(31 downto 0);  -- de2_pio_redled18_s1_translator:av_writedata -> de2_pio_redled18:writedata
	signal de2_pio_redled18_s1_translator_avalon_anti_slave_0_address                                                       : std_logic_vector(1 downto 0);   -- de2_pio_redled18_s1_translator:av_address -> de2_pio_redled18:address
	signal de2_pio_redled18_s1_translator_avalon_anti_slave_0_chipselect                                                    : std_logic;                      -- de2_pio_redled18_s1_translator:av_chipselect -> de2_pio_redled18:chipselect
	signal de2_pio_redled18_s1_translator_avalon_anti_slave_0_write                                                         : std_logic;                      -- de2_pio_redled18_s1_translator:av_write -> de2_pio_redled18_s1_translator_avalon_anti_slave_0_write:in
	signal de2_pio_redled18_s1_translator_avalon_anti_slave_0_readdata                                                      : std_logic_vector(31 downto 0);  -- de2_pio_redled18:readdata -> de2_pio_redled18_s1_translator:av_readdata
	signal de2_pio_greenled9_s1_translator_avalon_anti_slave_0_writedata                                                    : std_logic_vector(31 downto 0);  -- de2_pio_greenled9_s1_translator:av_writedata -> de2_pio_greenled9:writedata
	signal de2_pio_greenled9_s1_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(1 downto 0);   -- de2_pio_greenled9_s1_translator:av_address -> de2_pio_greenled9:address
	signal de2_pio_greenled9_s1_translator_avalon_anti_slave_0_chipselect                                                   : std_logic;                      -- de2_pio_greenled9_s1_translator:av_chipselect -> de2_pio_greenled9:chipselect
	signal de2_pio_greenled9_s1_translator_avalon_anti_slave_0_write                                                        : std_logic;                      -- de2_pio_greenled9_s1_translator:av_write -> de2_pio_greenled9_s1_translator_avalon_anti_slave_0_write:in
	signal de2_pio_greenled9_s1_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(31 downto 0);  -- de2_pio_greenled9:readdata -> de2_pio_greenled9_s1_translator:av_readdata
	signal de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_writedata                                                   : std_logic_vector(31 downto 0);  -- de2_pio_hex_high28_s1_translator:av_writedata -> de2_pio_hex_high28:writedata
	signal de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_address                                                     : std_logic_vector(1 downto 0);   -- de2_pio_hex_high28_s1_translator:av_address -> de2_pio_hex_high28:address
	signal de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_chipselect                                                  : std_logic;                      -- de2_pio_hex_high28_s1_translator:av_chipselect -> de2_pio_hex_high28:chipselect
	signal de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_write                                                       : std_logic;                      -- de2_pio_hex_high28_s1_translator:av_write -> de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_write:in
	signal de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_readdata                                                    : std_logic_vector(31 downto 0);  -- de2_pio_hex_high28:readdata -> de2_pio_hex_high28_s1_translator:av_readdata
	signal de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_writedata                                                    : std_logic_vector(31 downto 0);  -- de2_pio_hex_low28_s1_translator:av_writedata -> de2_pio_hex_low28:writedata
	signal de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(1 downto 0);   -- de2_pio_hex_low28_s1_translator:av_address -> de2_pio_hex_low28:address
	signal de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_chipselect                                                   : std_logic;                      -- de2_pio_hex_low28_s1_translator:av_chipselect -> de2_pio_hex_low28:chipselect
	signal de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_write                                                        : std_logic;                      -- de2_pio_hex_low28_s1_translator:av_write -> de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_write:in
	signal de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(31 downto 0);  -- de2_pio_hex_low28:readdata -> de2_pio_hex_low28_s1_translator:av_readdata
	signal sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata                                                  : std_logic_vector(15 downto 0);  -- sram_avalon_sram_slave_translator:av_writedata -> sram:writedata
	signal sram_avalon_sram_slave_translator_avalon_anti_slave_0_address                                                    : std_logic_vector(17 downto 0);  -- sram_avalon_sram_slave_translator:av_address -> sram:address
	signal sram_avalon_sram_slave_translator_avalon_anti_slave_0_write                                                      : std_logic;                      -- sram_avalon_sram_slave_translator:av_write -> sram:write
	signal sram_avalon_sram_slave_translator_avalon_anti_slave_0_read                                                       : std_logic;                      -- sram_avalon_sram_slave_translator:av_read -> sram:read
	signal sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata                                                   : std_logic_vector(15 downto 0);  -- sram:readdata -> sram_avalon_sram_slave_translator:av_readdata
	signal sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid                                              : std_logic;                      -- sram:readdatavalid -> sram_avalon_sram_slave_translator:av_readdatavalid
	signal sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable                                                 : std_logic_vector(1 downto 0);   -- sram_avalon_sram_slave_translator:av_byteenable -> sram:byteenable
	signal sdram_s1_translator_avalon_anti_slave_0_waitrequest                                                              : std_logic;                      -- sdram:za_waitrequest -> sdram_s1_translator:av_waitrequest
	signal sdram_s1_translator_avalon_anti_slave_0_writedata                                                                : std_logic_vector(15 downto 0);  -- sdram_s1_translator:av_writedata -> sdram:az_data
	signal sdram_s1_translator_avalon_anti_slave_0_address                                                                  : std_logic_vector(21 downto 0);  -- sdram_s1_translator:av_address -> sdram:az_addr
	signal sdram_s1_translator_avalon_anti_slave_0_chipselect                                                               : std_logic;                      -- sdram_s1_translator:av_chipselect -> sdram:az_cs
	signal sdram_s1_translator_avalon_anti_slave_0_write                                                                    : std_logic;                      -- sdram_s1_translator:av_write -> sdram_s1_translator_avalon_anti_slave_0_write:in
	signal sdram_s1_translator_avalon_anti_slave_0_read                                                                     : std_logic;                      -- sdram_s1_translator:av_read -> sdram_s1_translator_avalon_anti_slave_0_read:in
	signal sdram_s1_translator_avalon_anti_slave_0_readdata                                                                 : std_logic_vector(15 downto 0);  -- sdram:za_data -> sdram_s1_translator:av_readdata
	signal sdram_s1_translator_avalon_anti_slave_0_readdatavalid                                                            : std_logic;                      -- sdram:za_valid -> sdram_s1_translator:av_readdatavalid
	signal sdram_s1_translator_avalon_anti_slave_0_byteenable                                                               : std_logic_vector(1 downto 0);   -- sdram_s1_translator:av_byteenable -> sdram_s1_translator_avalon_anti_slave_0_byteenable:in
	signal nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_waitrequest                           : std_logic;                      -- nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_ht18_lemonde_streit_data_master_translator:uav_waitrequest
	signal nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_burstcount                            : std_logic_vector(2 downto 0);   -- nios2_ht18_lemonde_streit_data_master_translator:uav_burstcount -> nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_writedata                             : std_logic_vector(31 downto 0);  -- nios2_ht18_lemonde_streit_data_master_translator:uav_writedata -> nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_address                               : std_logic_vector(24 downto 0);  -- nios2_ht18_lemonde_streit_data_master_translator:uav_address -> nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:av_address
	signal nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_lock                                  : std_logic;                      -- nios2_ht18_lemonde_streit_data_master_translator:uav_lock -> nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_write                                 : std_logic;                      -- nios2_ht18_lemonde_streit_data_master_translator:uav_write -> nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:av_write
	signal nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_read                                  : std_logic;                      -- nios2_ht18_lemonde_streit_data_master_translator:uav_read -> nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:av_read
	signal nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_readdata                              : std_logic_vector(31 downto 0);  -- nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_ht18_lemonde_streit_data_master_translator:uav_readdata
	signal nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_debugaccess                           : std_logic;                      -- nios2_ht18_lemonde_streit_data_master_translator:uav_debugaccess -> nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_byteenable                            : std_logic_vector(3 downto 0);   -- nios2_ht18_lemonde_streit_data_master_translator:uav_byteenable -> nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_readdatavalid                         : std_logic;                      -- nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_ht18_lemonde_streit_data_master_translator:uav_readdatavalid
	signal nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_waitrequest                    : std_logic;                      -- nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_ht18_lemonde_streit_instruction_master_translator:uav_waitrequest
	signal nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_burstcount                     : std_logic_vector(2 downto 0);   -- nios2_ht18_lemonde_streit_instruction_master_translator:uav_burstcount -> nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_writedata                      : std_logic_vector(31 downto 0);  -- nios2_ht18_lemonde_streit_instruction_master_translator:uav_writedata -> nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_address                        : std_logic_vector(24 downto 0);  -- nios2_ht18_lemonde_streit_instruction_master_translator:uav_address -> nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_lock                           : std_logic;                      -- nios2_ht18_lemonde_streit_instruction_master_translator:uav_lock -> nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_write                          : std_logic;                      -- nios2_ht18_lemonde_streit_instruction_master_translator:uav_write -> nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_read                           : std_logic;                      -- nios2_ht18_lemonde_streit_instruction_master_translator:uav_read -> nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_readdata                       : std_logic_vector(31 downto 0);  -- nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_ht18_lemonde_streit_instruction_master_translator:uav_readdata
	signal nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_debugaccess                    : std_logic;                      -- nios2_ht18_lemonde_streit_instruction_master_translator:uav_debugaccess -> nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_byteenable                     : std_logic_vector(3 downto 0);   -- nios2_ht18_lemonde_streit_instruction_master_translator:uav_byteenable -> nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_readdatavalid                  : std_logic;                      -- nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_ht18_lemonde_streit_instruction_master_translator:uav_readdatavalid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                        : std_logic;                      -- onchip_memory_s1_translator:uav_waitrequest -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                         : std_logic_vector(2 downto 0);   -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory_s1_translator:uav_burstcount
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                          : std_logic_vector(31 downto 0);  -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory_s1_translator:uav_writedata
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address                                            : std_logic_vector(24 downto 0);  -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory_s1_translator:uav_address
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write                                              : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory_s1_translator:uav_write
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock                                               : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory_s1_translator:uav_lock
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read                                               : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory_s1_translator:uav_read
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                           : std_logic_vector(31 downto 0);  -- onchip_memory_s1_translator:uav_readdata -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                      : std_logic;                      -- onchip_memory_s1_translator:uav_readdatavalid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                        : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory_s1_translator:uav_debugaccess
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                         : std_logic_vector(3 downto 0);   -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory_s1_translator:uav_byteenable
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                 : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                       : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                               : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                        : std_logic_vector(100 downto 0); -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                       : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                              : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                    : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                            : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                     : std_logic_vector(100 downto 0); -- onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                    : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                  : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                   : std_logic_vector(33 downto 0);  -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                  : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                       : std_logic;                      -- ht18_lemonde_streit_control_slave_translator:uav_waitrequest -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                        : std_logic_vector(2 downto 0);   -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> ht18_lemonde_streit_control_slave_translator:uav_burstcount
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                         : std_logic_vector(31 downto 0);  -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> ht18_lemonde_streit_control_slave_translator:uav_writedata
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_address                           : std_logic_vector(24 downto 0);  -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> ht18_lemonde_streit_control_slave_translator:uav_address
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_write                             : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> ht18_lemonde_streit_control_slave_translator:uav_write
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                              : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> ht18_lemonde_streit_control_slave_translator:uav_lock
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_read                              : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> ht18_lemonde_streit_control_slave_translator:uav_read
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                          : std_logic_vector(31 downto 0);  -- ht18_lemonde_streit_control_slave_translator:uav_readdata -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                     : std_logic;                      -- ht18_lemonde_streit_control_slave_translator:uav_readdatavalid -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                       : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ht18_lemonde_streit_control_slave_translator:uav_debugaccess
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                        : std_logic_vector(3 downto 0);   -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> ht18_lemonde_streit_control_slave_translator:uav_byteenable
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                      : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket              : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                       : std_logic_vector(100 downto 0); -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                      : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket             : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                   : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket           : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                    : std_logic_vector(100 downto 0); -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                   : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                 : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                  : std_logic_vector(33 downto 0);  -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                 : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                           : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                            : std_logic_vector(2 downto 0);   -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata                             : std_logic_vector(31 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address                               : std_logic_vector(24 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write                                 : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock                                  : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read                                  : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata                              : std_logic_vector(31 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                         : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                           : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                            : std_logic_vector(3 downto 0);   -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                    : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                          : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                  : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data                           : std_logic_vector(100 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                          : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                 : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                       : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket               : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                        : std_logic_vector(100 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                       : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                     : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                      : std_logic_vector(33 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                     : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator:uav_waitrequest -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);   -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_ht18_lemonde_streit_jtag_debug_module_translator:uav_burstcount
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0);  -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_ht18_lemonde_streit_jtag_debug_module_translator:uav_writedata
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(24 downto 0);  -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_ht18_lemonde_streit_jtag_debug_module_translator:uav_address
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_ht18_lemonde_streit_jtag_debug_module_translator:uav_write
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_ht18_lemonde_streit_jtag_debug_module_translator:uav_lock
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_ht18_lemonde_streit_jtag_debug_module_translator:uav_read
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0);  -- nios2_ht18_lemonde_streit_jtag_debug_module_translator:uav_readdata -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator:uav_readdatavalid -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_ht18_lemonde_streit_jtag_debug_module_translator:uav_debugaccess
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);   -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_ht18_lemonde_streit_jtag_debug_module_translator:uav_byteenable
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(100 downto 0); -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(100 downto 0); -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0);  -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                              : std_logic;                      -- timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                               : std_logic_vector(2 downto 0);   -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                : std_logic_vector(31 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address                                                  : std_logic_vector(24 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write                                                    : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                     : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read                                                     : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                 : std_logic_vector(31 downto 0);  -- timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                            : std_logic;                      -- timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                              : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                               : std_logic_vector(3 downto 0);   -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                       : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                             : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                     : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                              : std_logic_vector(100 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                             : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                    : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                          : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                  : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                           : std_logic_vector(100 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                          : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                        : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                         : std_logic_vector(33 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                        : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                              : std_logic;                      -- timer_1_s1_translator:uav_waitrequest -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                               : std_logic_vector(2 downto 0);   -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_1_s1_translator:uav_burstcount
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                : std_logic_vector(31 downto 0);  -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_1_s1_translator:uav_writedata
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address                                                  : std_logic_vector(24 downto 0);  -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_1_s1_translator:uav_address
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write                                                    : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_1_s1_translator:uav_write
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                     : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_1_s1_translator:uav_lock
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read                                                     : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_1_s1_translator:uav_read
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                 : std_logic_vector(31 downto 0);  -- timer_1_s1_translator:uav_readdata -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                            : std_logic;                      -- timer_1_s1_translator:uav_readdatavalid -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                              : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_1_s1_translator:uav_debugaccess
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                               : std_logic_vector(3 downto 0);   -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_1_s1_translator:uav_byteenable
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                       : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                             : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                     : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                              : std_logic_vector(100 downto 0); -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                             : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                    : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                          : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                  : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                           : std_logic_vector(100 downto 0); -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                          : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                        : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                         : std_logic_vector(33 downto 0);  -- timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                        : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                      -- p_counter_control_slave_translator:uav_waitrequest -> p_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(2 downto 0);   -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> p_counter_control_slave_translator:uav_burstcount
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(31 downto 0);  -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> p_counter_control_slave_translator:uav_writedata
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(24 downto 0);  -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> p_counter_control_slave_translator:uav_address
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> p_counter_control_slave_translator:uav_write
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> p_counter_control_slave_translator:uav_lock
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> p_counter_control_slave_translator:uav_read
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(31 downto 0);  -- p_counter_control_slave_translator:uav_readdata -> p_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                      -- p_counter_control_slave_translator:uav_readdatavalid -> p_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> p_counter_control_slave_translator:uav_debugaccess
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(3 downto 0);   -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> p_counter_control_slave_translator:uav_byteenable
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(100 downto 0); -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> p_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> p_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> p_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> p_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(100 downto 0); -- p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> p_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> p_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(33 downto 0);  -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> p_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> p_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- de2_pio_toggles18_s1_translator:uav_waitrequest -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(2 downto 0);   -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> de2_pio_toggles18_s1_translator:uav_burstcount
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(31 downto 0);  -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> de2_pio_toggles18_s1_translator:uav_writedata
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:m0_address -> de2_pio_toggles18_s1_translator:uav_address
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:m0_write -> de2_pio_toggles18_s1_translator:uav_write
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:m0_lock -> de2_pio_toggles18_s1_translator:uav_lock
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:m0_read -> de2_pio_toggles18_s1_translator:uav_read
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(31 downto 0);  -- de2_pio_toggles18_s1_translator:uav_readdata -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- de2_pio_toggles18_s1_translator:uav_readdatavalid -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> de2_pio_toggles18_s1_translator:uav_debugaccess
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(3 downto 0);   -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> de2_pio_toggles18_s1_translator:uav_byteenable
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(100 downto 0); -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(100 downto 0); -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(33 downto 0);  -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                        : std_logic;                      -- de2_pio_keys4_s1_translator:uav_waitrequest -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                         : std_logic_vector(2 downto 0);   -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> de2_pio_keys4_s1_translator:uav_burstcount
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                          : std_logic_vector(31 downto 0);  -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> de2_pio_keys4_s1_translator:uav_writedata
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_address                                            : std_logic_vector(24 downto 0);  -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:m0_address -> de2_pio_keys4_s1_translator:uav_address
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_write                                              : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:m0_write -> de2_pio_keys4_s1_translator:uav_write
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_lock                                               : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:m0_lock -> de2_pio_keys4_s1_translator:uav_lock
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_read                                               : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:m0_read -> de2_pio_keys4_s1_translator:uav_read
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                           : std_logic_vector(31 downto 0);  -- de2_pio_keys4_s1_translator:uav_readdata -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                      : std_logic;                      -- de2_pio_keys4_s1_translator:uav_readdatavalid -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                        : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> de2_pio_keys4_s1_translator:uav_debugaccess
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                         : std_logic_vector(3 downto 0);   -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> de2_pio_keys4_s1_translator:uav_byteenable
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                 : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                       : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                               : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                        : std_logic_vector(100 downto 0); -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                       : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                              : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                    : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                            : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                     : std_logic_vector(100 downto 0); -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                    : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                  : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                   : std_logic_vector(33 downto 0);  -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                  : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                     : std_logic;                      -- de2_pio_redled18_s1_translator:uav_waitrequest -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                      : std_logic_vector(2 downto 0);   -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> de2_pio_redled18_s1_translator:uav_burstcount
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                       : std_logic_vector(31 downto 0);  -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> de2_pio_redled18_s1_translator:uav_writedata
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_address                                         : std_logic_vector(24 downto 0);  -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:m0_address -> de2_pio_redled18_s1_translator:uav_address
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_write                                           : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:m0_write -> de2_pio_redled18_s1_translator:uav_write
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_lock                                            : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:m0_lock -> de2_pio_redled18_s1_translator:uav_lock
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_read                                            : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:m0_read -> de2_pio_redled18_s1_translator:uav_read
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                        : std_logic_vector(31 downto 0);  -- de2_pio_redled18_s1_translator:uav_readdata -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                   : std_logic;                      -- de2_pio_redled18_s1_translator:uav_readdatavalid -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                     : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> de2_pio_redled18_s1_translator:uav_debugaccess
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                      : std_logic_vector(3 downto 0);   -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> de2_pio_redled18_s1_translator:uav_byteenable
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                              : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                    : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                            : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                     : std_logic_vector(100 downto 0); -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                    : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                           : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                 : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                         : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                  : std_logic_vector(100 downto 0); -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                 : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                               : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                : std_logic_vector(33 downto 0);  -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                               : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- de2_pio_greenled9_s1_translator:uav_waitrequest -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(2 downto 0);   -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> de2_pio_greenled9_s1_translator:uav_burstcount
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(31 downto 0);  -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> de2_pio_greenled9_s1_translator:uav_writedata
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:m0_address -> de2_pio_greenled9_s1_translator:uav_address
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:m0_write -> de2_pio_greenled9_s1_translator:uav_write
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:m0_lock -> de2_pio_greenled9_s1_translator:uav_lock
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:m0_read -> de2_pio_greenled9_s1_translator:uav_read
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(31 downto 0);  -- de2_pio_greenled9_s1_translator:uav_readdata -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- de2_pio_greenled9_s1_translator:uav_readdatavalid -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> de2_pio_greenled9_s1_translator:uav_debugaccess
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(3 downto 0);   -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> de2_pio_greenled9_s1_translator:uav_byteenable
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(100 downto 0); -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(100 downto 0); -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(33 downto 0);  -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                   : std_logic;                      -- de2_pio_hex_high28_s1_translator:uav_waitrequest -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                    : std_logic_vector(2 downto 0);   -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> de2_pio_hex_high28_s1_translator:uav_burstcount
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                     : std_logic_vector(31 downto 0);  -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> de2_pio_hex_high28_s1_translator:uav_writedata
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_address                                       : std_logic_vector(24 downto 0);  -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:m0_address -> de2_pio_hex_high28_s1_translator:uav_address
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_write                                         : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:m0_write -> de2_pio_hex_high28_s1_translator:uav_write
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_lock                                          : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:m0_lock -> de2_pio_hex_high28_s1_translator:uav_lock
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_read                                          : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:m0_read -> de2_pio_hex_high28_s1_translator:uav_read
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                      : std_logic_vector(31 downto 0);  -- de2_pio_hex_high28_s1_translator:uav_readdata -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                 : std_logic;                      -- de2_pio_hex_high28_s1_translator:uav_readdatavalid -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                   : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> de2_pio_hex_high28_s1_translator:uav_debugaccess
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                    : std_logic_vector(3 downto 0);   -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> de2_pio_hex_high28_s1_translator:uav_byteenable
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                            : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                  : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                          : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                   : std_logic_vector(100 downto 0); -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                  : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                         : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                               : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                       : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                : std_logic_vector(100 downto 0); -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                               : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                             : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                              : std_logic_vector(33 downto 0);  -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                             : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- de2_pio_hex_low28_s1_translator:uav_waitrequest -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(2 downto 0);   -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> de2_pio_hex_low28_s1_translator:uav_burstcount
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(31 downto 0);  -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> de2_pio_hex_low28_s1_translator:uav_writedata
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:m0_address -> de2_pio_hex_low28_s1_translator:uav_address
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:m0_write -> de2_pio_hex_low28_s1_translator:uav_write
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:m0_lock -> de2_pio_hex_low28_s1_translator:uav_lock
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:m0_read -> de2_pio_hex_low28_s1_translator:uav_read
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(31 downto 0);  -- de2_pio_hex_low28_s1_translator:uav_readdata -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- de2_pio_hex_low28_s1_translator:uav_readdatavalid -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> de2_pio_hex_low28_s1_translator:uav_debugaccess
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(3 downto 0);   -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> de2_pio_hex_low28_s1_translator:uav_byteenable
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(100 downto 0); -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(100 downto 0); -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(33 downto 0);  -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                                  : std_logic;                      -- sram_avalon_sram_slave_translator:uav_waitrequest -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                                   : std_logic_vector(1 downto 0);   -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sram_avalon_sram_slave_translator:uav_burstcount
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata                                    : std_logic_vector(15 downto 0);  -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sram_avalon_sram_slave_translator:uav_writedata
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address                                      : std_logic_vector(24 downto 0);  -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> sram_avalon_sram_slave_translator:uav_address
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write                                        : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> sram_avalon_sram_slave_translator:uav_write
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock                                         : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sram_avalon_sram_slave_translator:uav_lock
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read                                         : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> sram_avalon_sram_slave_translator:uav_read
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata                                     : std_logic_vector(15 downto 0);  -- sram_avalon_sram_slave_translator:uav_readdata -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                : std_logic;                      -- sram_avalon_sram_slave_translator:uav_readdatavalid -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                                  : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sram_avalon_sram_slave_translator:uav_debugaccess
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                                   : std_logic_vector(1 downto 0);   -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sram_avalon_sram_slave_translator:uav_byteenable
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                           : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                                 : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                         : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data                                  : std_logic_vector(82 downto 0);  -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                                 : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                        : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                              : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                      : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                               : std_logic_vector(82 downto 0);  -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                              : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                            : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                             : std_logic_vector(17 downto 0);  -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                            : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                            : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                             : std_logic_vector(17 downto 0);  -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                            : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                                : std_logic;                      -- sdram_s1_translator:uav_waitrequest -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                                 : std_logic_vector(1 downto 0);   -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_s1_translator:uav_burstcount
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                  : std_logic_vector(15 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_s1_translator:uav_writedata
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_address                                                    : std_logic_vector(24 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_s1_translator:uav_address
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_write                                                      : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_s1_translator:uav_write
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                       : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_s1_translator:uav_lock
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_read                                                       : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_s1_translator:uav_read
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                   : std_logic_vector(15 downto 0);  -- sdram_s1_translator:uav_readdata -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                              : std_logic;                      -- sdram_s1_translator:uav_readdatavalid -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                                : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_s1_translator:uav_debugaccess
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                                 : std_logic_vector(1 downto 0);   -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_s1_translator:uav_byteenable
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                         : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                               : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                       : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                                : std_logic_vector(82 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                               : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                      : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                            : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                    : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                             : std_logic_vector(82 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                            : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                          : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                           : std_logic_vector(17 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                          : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                                          : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                           : std_logic_vector(17 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                                          : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                  : std_logic;                      -- nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent_cp_valid                        : std_logic;                      -- nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                : std_logic;                      -- nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent_cp_data                         : std_logic_vector(99 downto 0);  -- nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent_cp_ready                        : std_logic;                      -- addr_router:sink_ready -> nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket           : std_logic;                      -- nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                 : std_logic;                      -- nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket         : std_logic;                      -- nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent_cp_data                  : std_logic_vector(99 downto 0);  -- nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                 : std_logic;                      -- addr_router_001:sink_ready -> nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                        : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid                                              : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                      : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data                                               : std_logic_vector(99 downto 0);  -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready                                              : std_logic;                      -- id_router:sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                       : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                             : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                     : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rp_data                              : std_logic_vector(99 downto 0);  -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                             : std_logic;                      -- id_router_001:sink_ready -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                           : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid                                 : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                         : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data                                  : std_logic_vector(99 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready                                 : std_logic;                      -- id_router_002:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(99 downto 0);  -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                      -- id_router_003:sink_ready -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                              : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                    : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                            : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data                                                     : std_logic_vector(99 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                    : std_logic;                      -- id_router_004:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                              : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                    : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                            : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data                                                     : std_logic_vector(99 downto 0);  -- timer_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                    : std_logic;                      -- id_router_005:sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(99 downto 0);  -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal p_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                      -- id_router_006:sink_ready -> p_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(99 downto 0);  -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	signal de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_007:sink_ready -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                        : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rp_valid                                              : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                      : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rp_data                                               : std_logic_vector(99 downto 0);  -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	signal de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rp_ready                                              : std_logic;                      -- id_router_008:sink_ready -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                     : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rp_valid                                           : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                   : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rp_data                                            : std_logic_vector(99 downto 0);  -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	signal de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rp_ready                                           : std_logic;                      -- id_router_009:sink_ready -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(99 downto 0);  -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	signal de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_010:sink_ready -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                   : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rp_valid                                         : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                 : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rp_data                                          : std_logic_vector(99 downto 0);  -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	signal de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rp_ready                                         : std_logic;                      -- id_router_011:sink_ready -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(99 downto 0);  -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	signal de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_012:sink_ready -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                                  : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid                                        : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                                : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data                                         : std_logic_vector(81 downto 0);  -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready                                        : std_logic;                      -- id_router_013:sink_ready -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                                : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                      : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                              : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_data                                                       : std_logic_vector(81 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                      : std_logic;                      -- id_router_014:sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal burst_adapter_source0_endofpacket                                                                                : std_logic;                      -- burst_adapter:source0_endofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_source0_valid                                                                                      : std_logic;                      -- burst_adapter:source0_valid -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_source0_startofpacket                                                                              : std_logic;                      -- burst_adapter:source0_startofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_source0_data                                                                                       : std_logic_vector(81 downto 0);  -- burst_adapter:source0_data -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_source0_ready                                                                                      : std_logic;                      -- sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	signal burst_adapter_source0_channel                                                                                    : std_logic_vector(14 downto 0);  -- burst_adapter:source0_channel -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_001_source0_endofpacket                                                                            : std_logic;                      -- burst_adapter_001:source0_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_001_source0_valid                                                                                  : std_logic;                      -- burst_adapter_001:source0_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_001_source0_startofpacket                                                                          : std_logic;                      -- burst_adapter_001:source0_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_001_source0_data                                                                                   : std_logic_vector(81 downto 0);  -- burst_adapter_001:source0_data -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_001_source0_ready                                                                                  : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	signal burst_adapter_001_source0_channel                                                                                : std_logic_vector(14 downto 0);  -- burst_adapter_001:source0_channel -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal rst_controller_reset_out_reset                                                                                   : std_logic;                      -- rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, burst_adapter:reset, burst_adapter_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_013:reset, cmd_xbar_mux_014:reset, de2_pio_greenled9_s1_translator:reset, de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:reset, de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, de2_pio_hex_high28_s1_translator:reset, de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:reset, de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, de2_pio_hex_low28_s1_translator:reset, de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:reset, de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, de2_pio_keys4_s1_translator:reset, de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:reset, de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, de2_pio_redled18_s1_translator:reset, de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:reset, de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, de2_pio_toggles18_s1_translator:reset, de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:reset, de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, irq_mapper:reset, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, nios2_ht18_lemonde_streit_data_master_translator:reset, nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:reset, nios2_ht18_lemonde_streit_instruction_master_translator:reset, nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_ht18_lemonde_streit_jtag_debug_module_translator:reset, nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory:reset, onchip_memory_s1_translator:reset, onchip_memory_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, p_counter_control_slave_translator:reset, p_counter_control_slave_translator_avalon_universal_slave_0_agent:reset, p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rst_controller_reset_out_reset:in, sdram_s1_translator:reset, sdram_s1_translator_avalon_universal_slave_0_agent:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sram:reset, sram_avalon_sram_slave_translator:reset, sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_1_s1_translator:reset, timer_1_s1_translator_avalon_universal_slave_0_agent:reset, timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset]
	signal rst_controller_reset_out_reset_req                                                                               : std_logic;                      -- rst_controller:reset_req -> onchip_memory:reset_req
	signal nios2_ht18_lemonde_streit_jtag_debug_module_reset_reset                                                          : std_logic;                      -- nios2_ht18_lemonde_streit:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller_002:reset_in1]
	signal rst_controller_001_reset_out_reset                                                                               : std_logic;                      -- rst_controller_001:reset_out -> [ht18_lemonde_streit_control_slave_translator:reset, ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:reset, ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_001:reset, rsp_xbar_demux_001:reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_002_reset_out_reset                                                                               : std_logic;                      -- rst_controller_002:reset_out -> up_clocks_0:reset
	signal cmd_xbar_demux_src0_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                                        : std_logic;                      -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                                      : std_logic_vector(14 downto 0);  -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                                        : std_logic;                      -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux:src1_endofpacket -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                                        : std_logic;                      -- cmd_xbar_demux:src1_valid -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux:src1_startofpacket -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_src1_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src1_data -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_src1_channel                                                                                      : std_logic_vector(14 downto 0);  -- cmd_xbar_demux:src1_channel -> ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_src2_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux:src2_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_src2_valid                                                                                        : std_logic;                      -- cmd_xbar_demux:src2_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_src2_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux:src2_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_src2_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src2_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_src2_channel                                                                                      : std_logic_vector(14 downto 0);  -- cmd_xbar_demux:src2_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_src3_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	signal cmd_xbar_demux_src3_valid                                                                                        : std_logic;                      -- cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	signal cmd_xbar_demux_src3_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	signal cmd_xbar_demux_src3_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	signal cmd_xbar_demux_src3_channel                                                                                      : std_logic_vector(14 downto 0);  -- cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	signal cmd_xbar_demux_src3_ready                                                                                        : std_logic;                      -- cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	signal cmd_xbar_demux_src4_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux:src4_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_src4_valid                                                                                        : std_logic;                      -- cmd_xbar_demux:src4_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_src4_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux:src4_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_src4_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src4_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_src4_channel                                                                                      : std_logic_vector(14 downto 0);  -- cmd_xbar_demux:src4_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_src5_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux:src5_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_src5_valid                                                                                        : std_logic;                      -- cmd_xbar_demux:src5_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_src5_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux:src5_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_src5_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src5_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_src5_channel                                                                                      : std_logic_vector(14 downto 0);  -- cmd_xbar_demux:src5_channel -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_src6_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux:src6_endofpacket -> p_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_src6_valid                                                                                        : std_logic;                      -- cmd_xbar_demux:src6_valid -> p_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_src6_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux:src6_startofpacket -> p_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_src6_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src6_data -> p_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_src6_channel                                                                                      : std_logic_vector(14 downto 0);  -- cmd_xbar_demux:src6_channel -> p_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_src7_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux:src7_endofpacket -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_src7_valid                                                                                        : std_logic;                      -- cmd_xbar_demux:src7_valid -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_src7_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux:src7_startofpacket -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_src7_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src7_data -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_src7_channel                                                                                      : std_logic_vector(14 downto 0);  -- cmd_xbar_demux:src7_channel -> de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_src8_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux:src8_endofpacket -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_src8_valid                                                                                        : std_logic;                      -- cmd_xbar_demux:src8_valid -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_src8_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux:src8_startofpacket -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_src8_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src8_data -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_src8_channel                                                                                      : std_logic_vector(14 downto 0);  -- cmd_xbar_demux:src8_channel -> de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_src9_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux:src9_endofpacket -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_src9_valid                                                                                        : std_logic;                      -- cmd_xbar_demux:src9_valid -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_src9_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux:src9_startofpacket -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_src9_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src9_data -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_src9_channel                                                                                      : std_logic_vector(14 downto 0);  -- cmd_xbar_demux:src9_channel -> de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_src10_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_demux:src10_endofpacket -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_src10_valid                                                                                       : std_logic;                      -- cmd_xbar_demux:src10_valid -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_src10_startofpacket                                                                               : std_logic;                      -- cmd_xbar_demux:src10_startofpacket -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_src10_data                                                                                        : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src10_data -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_src10_channel                                                                                     : std_logic_vector(14 downto 0);  -- cmd_xbar_demux:src10_channel -> de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_src11_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_demux:src11_endofpacket -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_src11_valid                                                                                       : std_logic;                      -- cmd_xbar_demux:src11_valid -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_src11_startofpacket                                                                               : std_logic;                      -- cmd_xbar_demux:src11_startofpacket -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_src11_data                                                                                        : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src11_data -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_src11_channel                                                                                     : std_logic_vector(14 downto 0);  -- cmd_xbar_demux:src11_channel -> de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_src12_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_demux:src12_endofpacket -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_src12_valid                                                                                       : std_logic;                      -- cmd_xbar_demux:src12_valid -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_src12_startofpacket                                                                               : std_logic;                      -- cmd_xbar_demux:src12_startofpacket -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_src12_data                                                                                        : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src12_data -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_src12_channel                                                                                     : std_logic_vector(14 downto 0);  -- cmd_xbar_demux:src12_channel -> de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_src13_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_demux:src13_endofpacket -> cmd_xbar_mux_013:sink0_endofpacket
	signal cmd_xbar_demux_src13_valid                                                                                       : std_logic;                      -- cmd_xbar_demux:src13_valid -> cmd_xbar_mux_013:sink0_valid
	signal cmd_xbar_demux_src13_startofpacket                                                                               : std_logic;                      -- cmd_xbar_demux:src13_startofpacket -> cmd_xbar_mux_013:sink0_startofpacket
	signal cmd_xbar_demux_src13_data                                                                                        : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src13_data -> cmd_xbar_mux_013:sink0_data
	signal cmd_xbar_demux_src13_channel                                                                                     : std_logic_vector(14 downto 0);  -- cmd_xbar_demux:src13_channel -> cmd_xbar_mux_013:sink0_channel
	signal cmd_xbar_demux_src13_ready                                                                                       : std_logic;                      -- cmd_xbar_mux_013:sink0_ready -> cmd_xbar_demux:src13_ready
	signal cmd_xbar_demux_src14_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_demux:src14_endofpacket -> cmd_xbar_mux_014:sink0_endofpacket
	signal cmd_xbar_demux_src14_valid                                                                                       : std_logic;                      -- cmd_xbar_demux:src14_valid -> cmd_xbar_mux_014:sink0_valid
	signal cmd_xbar_demux_src14_startofpacket                                                                               : std_logic;                      -- cmd_xbar_demux:src14_startofpacket -> cmd_xbar_mux_014:sink0_startofpacket
	signal cmd_xbar_demux_src14_data                                                                                        : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src14_data -> cmd_xbar_mux_014:sink0_data
	signal cmd_xbar_demux_src14_channel                                                                                     : std_logic_vector(14 downto 0);  -- cmd_xbar_demux:src14_channel -> cmd_xbar_mux_014:sink0_channel
	signal cmd_xbar_demux_src14_ready                                                                                       : std_logic;                      -- cmd_xbar_mux_014:sink0_ready -> cmd_xbar_demux:src14_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                                              : std_logic;                      -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                                    : std_logic;                      -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                                            : std_logic;                      -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                                     : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                                                  : std_logic_vector(14 downto 0);  -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                                    : std_logic;                      -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                                              : std_logic;                      -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                                                    : std_logic;                      -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_003:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                                            : std_logic;                      -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                                                     : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_003:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                                                  : std_logic_vector(14 downto 0);  -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_003:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                                                    : std_logic;                      -- cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal cmd_xbar_demux_001_src2_endofpacket                                                                              : std_logic;                      -- cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_013:sink1_endofpacket
	signal cmd_xbar_demux_001_src2_valid                                                                                    : std_logic;                      -- cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_013:sink1_valid
	signal cmd_xbar_demux_001_src2_startofpacket                                                                            : std_logic;                      -- cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_013:sink1_startofpacket
	signal cmd_xbar_demux_001_src2_data                                                                                     : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_013:sink1_data
	signal cmd_xbar_demux_001_src2_channel                                                                                  : std_logic_vector(14 downto 0);  -- cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_013:sink1_channel
	signal cmd_xbar_demux_001_src2_ready                                                                                    : std_logic;                      -- cmd_xbar_mux_013:sink1_ready -> cmd_xbar_demux_001:src2_ready
	signal cmd_xbar_demux_001_src3_endofpacket                                                                              : std_logic;                      -- cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_014:sink1_endofpacket
	signal cmd_xbar_demux_001_src3_valid                                                                                    : std_logic;                      -- cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_014:sink1_valid
	signal cmd_xbar_demux_001_src3_startofpacket                                                                            : std_logic;                      -- cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_014:sink1_startofpacket
	signal cmd_xbar_demux_001_src3_data                                                                                     : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_014:sink1_data
	signal cmd_xbar_demux_001_src3_channel                                                                                  : std_logic_vector(14 downto 0);  -- cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_014:sink1_channel
	signal cmd_xbar_demux_001_src3_ready                                                                                    : std_logic;                      -- cmd_xbar_mux_014:sink1_ready -> cmd_xbar_demux_001:src3_ready
	signal rsp_xbar_demux_src0_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                                        : std_logic;                      -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                                      : std_logic_vector(14 downto 0);  -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                                        : std_logic;                      -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                                        : std_logic;                      -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                                      : std_logic_vector(14 downto 0);  -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                                        : std_logic;                      -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                                              : std_logic;                      -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                                    : std_logic;                      -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                                            : std_logic;                      -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                                     : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                                                  : std_logic_vector(14 downto 0);  -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                                    : std_logic;                      -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_002_src0_endofpacket                                                                              : std_logic;                      -- rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                                    : std_logic;                      -- rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                                            : std_logic;                      -- rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                                     : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	signal rsp_xbar_demux_002_src0_channel                                                                                  : std_logic_vector(14 downto 0);  -- rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	signal rsp_xbar_demux_002_src0_ready                                                                                    : std_logic;                      -- rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	signal rsp_xbar_demux_003_src0_endofpacket                                                                              : std_logic;                      -- rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                                    : std_logic;                      -- rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                                            : std_logic;                      -- rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                                     : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	signal rsp_xbar_demux_003_src0_channel                                                                                  : std_logic_vector(14 downto 0);  -- rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	signal rsp_xbar_demux_003_src0_ready                                                                                    : std_logic;                      -- rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	signal rsp_xbar_demux_003_src1_endofpacket                                                                              : std_logic;                      -- rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_003_src1_valid                                                                                    : std_logic;                      -- rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_003_src1_startofpacket                                                                            : std_logic;                      -- rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_003_src1_data                                                                                     : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_003_src1_channel                                                                                  : std_logic_vector(14 downto 0);  -- rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_003_src1_ready                                                                                    : std_logic;                      -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_003:src1_ready
	signal rsp_xbar_demux_004_src0_endofpacket                                                                              : std_logic;                      -- rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                                    : std_logic;                      -- rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                                            : std_logic;                      -- rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                                     : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	signal rsp_xbar_demux_004_src0_channel                                                                                  : std_logic_vector(14 downto 0);  -- rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	signal rsp_xbar_demux_004_src0_ready                                                                                    : std_logic;                      -- rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	signal rsp_xbar_demux_005_src0_endofpacket                                                                              : std_logic;                      -- rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                                    : std_logic;                      -- rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                                            : std_logic;                      -- rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                                     : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	signal rsp_xbar_demux_005_src0_channel                                                                                  : std_logic_vector(14 downto 0);  -- rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	signal rsp_xbar_demux_005_src0_ready                                                                                    : std_logic;                      -- rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	signal rsp_xbar_demux_006_src0_endofpacket                                                                              : std_logic;                      -- rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                                    : std_logic;                      -- rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                                            : std_logic;                      -- rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                                     : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	signal rsp_xbar_demux_006_src0_channel                                                                                  : std_logic_vector(14 downto 0);  -- rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	signal rsp_xbar_demux_006_src0_ready                                                                                    : std_logic;                      -- rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	signal rsp_xbar_demux_007_src0_endofpacket                                                                              : std_logic;                      -- rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux:sink7_endofpacket
	signal rsp_xbar_demux_007_src0_valid                                                                                    : std_logic;                      -- rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux:sink7_valid
	signal rsp_xbar_demux_007_src0_startofpacket                                                                            : std_logic;                      -- rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux:sink7_startofpacket
	signal rsp_xbar_demux_007_src0_data                                                                                     : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_007:src0_data -> rsp_xbar_mux:sink7_data
	signal rsp_xbar_demux_007_src0_channel                                                                                  : std_logic_vector(14 downto 0);  -- rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux:sink7_channel
	signal rsp_xbar_demux_007_src0_ready                                                                                    : std_logic;                      -- rsp_xbar_mux:sink7_ready -> rsp_xbar_demux_007:src0_ready
	signal rsp_xbar_demux_008_src0_endofpacket                                                                              : std_logic;                      -- rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux:sink8_endofpacket
	signal rsp_xbar_demux_008_src0_valid                                                                                    : std_logic;                      -- rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux:sink8_valid
	signal rsp_xbar_demux_008_src0_startofpacket                                                                            : std_logic;                      -- rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux:sink8_startofpacket
	signal rsp_xbar_demux_008_src0_data                                                                                     : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_008:src0_data -> rsp_xbar_mux:sink8_data
	signal rsp_xbar_demux_008_src0_channel                                                                                  : std_logic_vector(14 downto 0);  -- rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux:sink8_channel
	signal rsp_xbar_demux_008_src0_ready                                                                                    : std_logic;                      -- rsp_xbar_mux:sink8_ready -> rsp_xbar_demux_008:src0_ready
	signal rsp_xbar_demux_009_src0_endofpacket                                                                              : std_logic;                      -- rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux:sink9_endofpacket
	signal rsp_xbar_demux_009_src0_valid                                                                                    : std_logic;                      -- rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux:sink9_valid
	signal rsp_xbar_demux_009_src0_startofpacket                                                                            : std_logic;                      -- rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux:sink9_startofpacket
	signal rsp_xbar_demux_009_src0_data                                                                                     : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_009:src0_data -> rsp_xbar_mux:sink9_data
	signal rsp_xbar_demux_009_src0_channel                                                                                  : std_logic_vector(14 downto 0);  -- rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux:sink9_channel
	signal rsp_xbar_demux_009_src0_ready                                                                                    : std_logic;                      -- rsp_xbar_mux:sink9_ready -> rsp_xbar_demux_009:src0_ready
	signal rsp_xbar_demux_010_src0_endofpacket                                                                              : std_logic;                      -- rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux:sink10_endofpacket
	signal rsp_xbar_demux_010_src0_valid                                                                                    : std_logic;                      -- rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux:sink10_valid
	signal rsp_xbar_demux_010_src0_startofpacket                                                                            : std_logic;                      -- rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux:sink10_startofpacket
	signal rsp_xbar_demux_010_src0_data                                                                                     : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_010:src0_data -> rsp_xbar_mux:sink10_data
	signal rsp_xbar_demux_010_src0_channel                                                                                  : std_logic_vector(14 downto 0);  -- rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux:sink10_channel
	signal rsp_xbar_demux_010_src0_ready                                                                                    : std_logic;                      -- rsp_xbar_mux:sink10_ready -> rsp_xbar_demux_010:src0_ready
	signal rsp_xbar_demux_011_src0_endofpacket                                                                              : std_logic;                      -- rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux:sink11_endofpacket
	signal rsp_xbar_demux_011_src0_valid                                                                                    : std_logic;                      -- rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux:sink11_valid
	signal rsp_xbar_demux_011_src0_startofpacket                                                                            : std_logic;                      -- rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux:sink11_startofpacket
	signal rsp_xbar_demux_011_src0_data                                                                                     : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_011:src0_data -> rsp_xbar_mux:sink11_data
	signal rsp_xbar_demux_011_src0_channel                                                                                  : std_logic_vector(14 downto 0);  -- rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux:sink11_channel
	signal rsp_xbar_demux_011_src0_ready                                                                                    : std_logic;                      -- rsp_xbar_mux:sink11_ready -> rsp_xbar_demux_011:src0_ready
	signal rsp_xbar_demux_012_src0_endofpacket                                                                              : std_logic;                      -- rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux:sink12_endofpacket
	signal rsp_xbar_demux_012_src0_valid                                                                                    : std_logic;                      -- rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux:sink12_valid
	signal rsp_xbar_demux_012_src0_startofpacket                                                                            : std_logic;                      -- rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux:sink12_startofpacket
	signal rsp_xbar_demux_012_src0_data                                                                                     : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_012:src0_data -> rsp_xbar_mux:sink12_data
	signal rsp_xbar_demux_012_src0_channel                                                                                  : std_logic_vector(14 downto 0);  -- rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux:sink12_channel
	signal rsp_xbar_demux_012_src0_ready                                                                                    : std_logic;                      -- rsp_xbar_mux:sink12_ready -> rsp_xbar_demux_012:src0_ready
	signal rsp_xbar_demux_013_src0_endofpacket                                                                              : std_logic;                      -- rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux:sink13_endofpacket
	signal rsp_xbar_demux_013_src0_valid                                                                                    : std_logic;                      -- rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux:sink13_valid
	signal rsp_xbar_demux_013_src0_startofpacket                                                                            : std_logic;                      -- rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux:sink13_startofpacket
	signal rsp_xbar_demux_013_src0_data                                                                                     : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_013:src0_data -> rsp_xbar_mux:sink13_data
	signal rsp_xbar_demux_013_src0_channel                                                                                  : std_logic_vector(14 downto 0);  -- rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux:sink13_channel
	signal rsp_xbar_demux_013_src0_ready                                                                                    : std_logic;                      -- rsp_xbar_mux:sink13_ready -> rsp_xbar_demux_013:src0_ready
	signal rsp_xbar_demux_013_src1_endofpacket                                                                              : std_logic;                      -- rsp_xbar_demux_013:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	signal rsp_xbar_demux_013_src1_valid                                                                                    : std_logic;                      -- rsp_xbar_demux_013:src1_valid -> rsp_xbar_mux_001:sink2_valid
	signal rsp_xbar_demux_013_src1_startofpacket                                                                            : std_logic;                      -- rsp_xbar_demux_013:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	signal rsp_xbar_demux_013_src1_data                                                                                     : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_013:src1_data -> rsp_xbar_mux_001:sink2_data
	signal rsp_xbar_demux_013_src1_channel                                                                                  : std_logic_vector(14 downto 0);  -- rsp_xbar_demux_013:src1_channel -> rsp_xbar_mux_001:sink2_channel
	signal rsp_xbar_demux_013_src1_ready                                                                                    : std_logic;                      -- rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_013:src1_ready
	signal rsp_xbar_demux_014_src0_endofpacket                                                                              : std_logic;                      -- rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux:sink14_endofpacket
	signal rsp_xbar_demux_014_src0_valid                                                                                    : std_logic;                      -- rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux:sink14_valid
	signal rsp_xbar_demux_014_src0_startofpacket                                                                            : std_logic;                      -- rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux:sink14_startofpacket
	signal rsp_xbar_demux_014_src0_data                                                                                     : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_014:src0_data -> rsp_xbar_mux:sink14_data
	signal rsp_xbar_demux_014_src0_channel                                                                                  : std_logic_vector(14 downto 0);  -- rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux:sink14_channel
	signal rsp_xbar_demux_014_src0_ready                                                                                    : std_logic;                      -- rsp_xbar_mux:sink14_ready -> rsp_xbar_demux_014:src0_ready
	signal rsp_xbar_demux_014_src1_endofpacket                                                                              : std_logic;                      -- rsp_xbar_demux_014:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	signal rsp_xbar_demux_014_src1_valid                                                                                    : std_logic;                      -- rsp_xbar_demux_014:src1_valid -> rsp_xbar_mux_001:sink3_valid
	signal rsp_xbar_demux_014_src1_startofpacket                                                                            : std_logic;                      -- rsp_xbar_demux_014:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	signal rsp_xbar_demux_014_src1_data                                                                                     : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_014:src1_data -> rsp_xbar_mux_001:sink3_data
	signal rsp_xbar_demux_014_src1_channel                                                                                  : std_logic_vector(14 downto 0);  -- rsp_xbar_demux_014:src1_channel -> rsp_xbar_mux_001:sink3_channel
	signal rsp_xbar_demux_014_src1_ready                                                                                    : std_logic;                      -- rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_014:src1_ready
	signal addr_router_src_endofpacket                                                                                      : std_logic;                      -- addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal addr_router_src_valid                                                                                            : std_logic;                      -- addr_router:src_valid -> cmd_xbar_demux:sink_valid
	signal addr_router_src_startofpacket                                                                                    : std_logic;                      -- addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal addr_router_src_data                                                                                             : std_logic_vector(99 downto 0);  -- addr_router:src_data -> cmd_xbar_demux:sink_data
	signal addr_router_src_channel                                                                                          : std_logic_vector(14 downto 0);  -- addr_router:src_channel -> cmd_xbar_demux:sink_channel
	signal addr_router_src_ready                                                                                            : std_logic;                      -- cmd_xbar_demux:sink_ready -> addr_router:src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                                     : std_logic;                      -- rsp_xbar_mux:src_endofpacket -> nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_src_valid                                                                                           : std_logic;                      -- rsp_xbar_mux:src_valid -> nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_src_startofpacket                                                                                   : std_logic;                      -- rsp_xbar_mux:src_startofpacket -> nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_src_data                                                                                            : std_logic_vector(99 downto 0);  -- rsp_xbar_mux:src_data -> nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_src_channel                                                                                         : std_logic_vector(14 downto 0);  -- rsp_xbar_mux:src_channel -> nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_src_ready                                                                                           : std_logic;                      -- nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	signal addr_router_001_src_endofpacket                                                                                  : std_logic;                      -- addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal addr_router_001_src_valid                                                                                        : std_logic;                      -- addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	signal addr_router_001_src_startofpacket                                                                                : std_logic;                      -- addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal addr_router_001_src_data                                                                                         : std_logic_vector(99 downto 0);  -- addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	signal addr_router_001_src_channel                                                                                      : std_logic_vector(14 downto 0);  -- addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	signal addr_router_001_src_ready                                                                                        : std_logic;                      -- cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_mux_001:src_endofpacket -> nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                                       : std_logic;                      -- rsp_xbar_mux_001:src_valid -> nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                                               : std_logic;                      -- rsp_xbar_mux_001:src_startofpacket -> nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                                        : std_logic_vector(99 downto 0);  -- rsp_xbar_mux_001:src_data -> nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_001_src_channel                                                                                     : std_logic_vector(14 downto 0);  -- rsp_xbar_mux_001:src_channel -> nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_001_src_ready                                                                                       : std_logic;                      -- nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	signal cmd_xbar_mux_src_endofpacket                                                                                     : std_logic;                      -- cmd_xbar_mux:src_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_src_valid                                                                                           : std_logic;                      -- cmd_xbar_mux:src_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_src_startofpacket                                                                                   : std_logic;                      -- cmd_xbar_mux:src_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_src_data                                                                                            : std_logic_vector(99 downto 0);  -- cmd_xbar_mux:src_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_src_channel                                                                                         : std_logic_vector(14 downto 0);  -- cmd_xbar_mux:src_channel -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_src_ready                                                                                           : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                                        : std_logic;                      -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                                              : std_logic;                      -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                                      : std_logic;                      -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                                               : std_logic_vector(99 downto 0);  -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                                            : std_logic_vector(14 downto 0);  -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                                              : std_logic;                      -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_demux_src1_ready                                                                                        : std_logic;                      -- ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src1_ready
	signal id_router_001_src_endofpacket                                                                                    : std_logic;                      -- id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal id_router_001_src_valid                                                                                          : std_logic;                      -- id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	signal id_router_001_src_startofpacket                                                                                  : std_logic;                      -- id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal id_router_001_src_data                                                                                           : std_logic_vector(99 downto 0);  -- id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	signal id_router_001_src_channel                                                                                        : std_logic_vector(14 downto 0);  -- id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	signal id_router_001_src_ready                                                                                          : std_logic;                      -- rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	signal cmd_xbar_demux_src2_ready                                                                                        : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src2_ready
	signal id_router_002_src_endofpacket                                                                                    : std_logic;                      -- id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal id_router_002_src_valid                                                                                          : std_logic;                      -- id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	signal id_router_002_src_startofpacket                                                                                  : std_logic;                      -- id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal id_router_002_src_data                                                                                           : std_logic_vector(99 downto 0);  -- id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	signal id_router_002_src_channel                                                                                        : std_logic_vector(14 downto 0);  -- id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	signal id_router_002_src_ready                                                                                          : std_logic;                      -- rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	signal cmd_xbar_mux_003_src_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_mux_003:src_endofpacket -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_003_src_valid                                                                                       : std_logic;                      -- cmd_xbar_mux_003:src_valid -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_003_src_startofpacket                                                                               : std_logic;                      -- cmd_xbar_mux_003:src_startofpacket -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_003_src_data                                                                                        : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_003:src_data -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_003_src_channel                                                                                     : std_logic_vector(14 downto 0);  -- cmd_xbar_mux_003:src_channel -> nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_003_src_ready                                                                                       : std_logic;                      -- nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	signal id_router_003_src_endofpacket                                                                                    : std_logic;                      -- id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal id_router_003_src_valid                                                                                          : std_logic;                      -- id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	signal id_router_003_src_startofpacket                                                                                  : std_logic;                      -- id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal id_router_003_src_data                                                                                           : std_logic_vector(99 downto 0);  -- id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	signal id_router_003_src_channel                                                                                        : std_logic_vector(14 downto 0);  -- id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	signal id_router_003_src_ready                                                                                          : std_logic;                      -- rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	signal cmd_xbar_demux_src4_ready                                                                                        : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src4_ready
	signal id_router_004_src_endofpacket                                                                                    : std_logic;                      -- id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal id_router_004_src_valid                                                                                          : std_logic;                      -- id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	signal id_router_004_src_startofpacket                                                                                  : std_logic;                      -- id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal id_router_004_src_data                                                                                           : std_logic_vector(99 downto 0);  -- id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	signal id_router_004_src_channel                                                                                        : std_logic_vector(14 downto 0);  -- id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	signal id_router_004_src_ready                                                                                          : std_logic;                      -- rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	signal cmd_xbar_demux_src5_ready                                                                                        : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src5_ready
	signal id_router_005_src_endofpacket                                                                                    : std_logic;                      -- id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal id_router_005_src_valid                                                                                          : std_logic;                      -- id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	signal id_router_005_src_startofpacket                                                                                  : std_logic;                      -- id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal id_router_005_src_data                                                                                           : std_logic_vector(99 downto 0);  -- id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	signal id_router_005_src_channel                                                                                        : std_logic_vector(14 downto 0);  -- id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	signal id_router_005_src_ready                                                                                          : std_logic;                      -- rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	signal cmd_xbar_demux_src6_ready                                                                                        : std_logic;                      -- p_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src6_ready
	signal id_router_006_src_endofpacket                                                                                    : std_logic;                      -- id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal id_router_006_src_valid                                                                                          : std_logic;                      -- id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	signal id_router_006_src_startofpacket                                                                                  : std_logic;                      -- id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal id_router_006_src_data                                                                                           : std_logic_vector(99 downto 0);  -- id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	signal id_router_006_src_channel                                                                                        : std_logic_vector(14 downto 0);  -- id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	signal id_router_006_src_ready                                                                                          : std_logic;                      -- rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	signal cmd_xbar_demux_src7_ready                                                                                        : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src7_ready
	signal id_router_007_src_endofpacket                                                                                    : std_logic;                      -- id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	signal id_router_007_src_valid                                                                                          : std_logic;                      -- id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	signal id_router_007_src_startofpacket                                                                                  : std_logic;                      -- id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	signal id_router_007_src_data                                                                                           : std_logic_vector(99 downto 0);  -- id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	signal id_router_007_src_channel                                                                                        : std_logic_vector(14 downto 0);  -- id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	signal id_router_007_src_ready                                                                                          : std_logic;                      -- rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	signal cmd_xbar_demux_src8_ready                                                                                        : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src8_ready
	signal id_router_008_src_endofpacket                                                                                    : std_logic;                      -- id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	signal id_router_008_src_valid                                                                                          : std_logic;                      -- id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	signal id_router_008_src_startofpacket                                                                                  : std_logic;                      -- id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	signal id_router_008_src_data                                                                                           : std_logic_vector(99 downto 0);  -- id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	signal id_router_008_src_channel                                                                                        : std_logic_vector(14 downto 0);  -- id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	signal id_router_008_src_ready                                                                                          : std_logic;                      -- rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	signal cmd_xbar_demux_src9_ready                                                                                        : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src9_ready
	signal id_router_009_src_endofpacket                                                                                    : std_logic;                      -- id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	signal id_router_009_src_valid                                                                                          : std_logic;                      -- id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	signal id_router_009_src_startofpacket                                                                                  : std_logic;                      -- id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	signal id_router_009_src_data                                                                                           : std_logic_vector(99 downto 0);  -- id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	signal id_router_009_src_channel                                                                                        : std_logic_vector(14 downto 0);  -- id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	signal id_router_009_src_ready                                                                                          : std_logic;                      -- rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	signal cmd_xbar_demux_src10_ready                                                                                       : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src10_ready
	signal id_router_010_src_endofpacket                                                                                    : std_logic;                      -- id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	signal id_router_010_src_valid                                                                                          : std_logic;                      -- id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	signal id_router_010_src_startofpacket                                                                                  : std_logic;                      -- id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	signal id_router_010_src_data                                                                                           : std_logic_vector(99 downto 0);  -- id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	signal id_router_010_src_channel                                                                                        : std_logic_vector(14 downto 0);  -- id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	signal id_router_010_src_ready                                                                                          : std_logic;                      -- rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	signal cmd_xbar_demux_src11_ready                                                                                       : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src11_ready
	signal id_router_011_src_endofpacket                                                                                    : std_logic;                      -- id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	signal id_router_011_src_valid                                                                                          : std_logic;                      -- id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	signal id_router_011_src_startofpacket                                                                                  : std_logic;                      -- id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	signal id_router_011_src_data                                                                                           : std_logic_vector(99 downto 0);  -- id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	signal id_router_011_src_channel                                                                                        : std_logic_vector(14 downto 0);  -- id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	signal id_router_011_src_ready                                                                                          : std_logic;                      -- rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	signal cmd_xbar_demux_src12_ready                                                                                       : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src12_ready
	signal id_router_012_src_endofpacket                                                                                    : std_logic;                      -- id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	signal id_router_012_src_valid                                                                                          : std_logic;                      -- id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	signal id_router_012_src_startofpacket                                                                                  : std_logic;                      -- id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	signal id_router_012_src_data                                                                                           : std_logic_vector(99 downto 0);  -- id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	signal id_router_012_src_channel                                                                                        : std_logic_vector(14 downto 0);  -- id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	signal id_router_012_src_ready                                                                                          : std_logic;                      -- rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	signal cmd_xbar_mux_013_src_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_mux_013:src_endofpacket -> width_adapter:in_endofpacket
	signal cmd_xbar_mux_013_src_valid                                                                                       : std_logic;                      -- cmd_xbar_mux_013:src_valid -> width_adapter:in_valid
	signal cmd_xbar_mux_013_src_startofpacket                                                                               : std_logic;                      -- cmd_xbar_mux_013:src_startofpacket -> width_adapter:in_startofpacket
	signal cmd_xbar_mux_013_src_data                                                                                        : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_013:src_data -> width_adapter:in_data
	signal cmd_xbar_mux_013_src_channel                                                                                     : std_logic_vector(14 downto 0);  -- cmd_xbar_mux_013:src_channel -> width_adapter:in_channel
	signal cmd_xbar_mux_013_src_ready                                                                                       : std_logic;                      -- width_adapter:in_ready -> cmd_xbar_mux_013:src_ready
	signal width_adapter_src_endofpacket                                                                                    : std_logic;                      -- width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	signal width_adapter_src_valid                                                                                          : std_logic;                      -- width_adapter:out_valid -> burst_adapter:sink0_valid
	signal width_adapter_src_startofpacket                                                                                  : std_logic;                      -- width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	signal width_adapter_src_data                                                                                           : std_logic_vector(81 downto 0);  -- width_adapter:out_data -> burst_adapter:sink0_data
	signal width_adapter_src_ready                                                                                          : std_logic;                      -- burst_adapter:sink0_ready -> width_adapter:out_ready
	signal width_adapter_src_channel                                                                                        : std_logic_vector(14 downto 0);  -- width_adapter:out_channel -> burst_adapter:sink0_channel
	signal id_router_013_src_endofpacket                                                                                    : std_logic;                      -- id_router_013:src_endofpacket -> width_adapter_001:in_endofpacket
	signal id_router_013_src_valid                                                                                          : std_logic;                      -- id_router_013:src_valid -> width_adapter_001:in_valid
	signal id_router_013_src_startofpacket                                                                                  : std_logic;                      -- id_router_013:src_startofpacket -> width_adapter_001:in_startofpacket
	signal id_router_013_src_data                                                                                           : std_logic_vector(81 downto 0);  -- id_router_013:src_data -> width_adapter_001:in_data
	signal id_router_013_src_channel                                                                                        : std_logic_vector(14 downto 0);  -- id_router_013:src_channel -> width_adapter_001:in_channel
	signal id_router_013_src_ready                                                                                          : std_logic;                      -- width_adapter_001:in_ready -> id_router_013:src_ready
	signal width_adapter_001_src_endofpacket                                                                                : std_logic;                      -- width_adapter_001:out_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	signal width_adapter_001_src_valid                                                                                      : std_logic;                      -- width_adapter_001:out_valid -> rsp_xbar_demux_013:sink_valid
	signal width_adapter_001_src_startofpacket                                                                              : std_logic;                      -- width_adapter_001:out_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	signal width_adapter_001_src_data                                                                                       : std_logic_vector(99 downto 0);  -- width_adapter_001:out_data -> rsp_xbar_demux_013:sink_data
	signal width_adapter_001_src_ready                                                                                      : std_logic;                      -- rsp_xbar_demux_013:sink_ready -> width_adapter_001:out_ready
	signal width_adapter_001_src_channel                                                                                    : std_logic_vector(14 downto 0);  -- width_adapter_001:out_channel -> rsp_xbar_demux_013:sink_channel
	signal cmd_xbar_mux_014_src_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_mux_014:src_endofpacket -> width_adapter_002:in_endofpacket
	signal cmd_xbar_mux_014_src_valid                                                                                       : std_logic;                      -- cmd_xbar_mux_014:src_valid -> width_adapter_002:in_valid
	signal cmd_xbar_mux_014_src_startofpacket                                                                               : std_logic;                      -- cmd_xbar_mux_014:src_startofpacket -> width_adapter_002:in_startofpacket
	signal cmd_xbar_mux_014_src_data                                                                                        : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_014:src_data -> width_adapter_002:in_data
	signal cmd_xbar_mux_014_src_channel                                                                                     : std_logic_vector(14 downto 0);  -- cmd_xbar_mux_014:src_channel -> width_adapter_002:in_channel
	signal cmd_xbar_mux_014_src_ready                                                                                       : std_logic;                      -- width_adapter_002:in_ready -> cmd_xbar_mux_014:src_ready
	signal width_adapter_002_src_endofpacket                                                                                : std_logic;                      -- width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	signal width_adapter_002_src_valid                                                                                      : std_logic;                      -- width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	signal width_adapter_002_src_startofpacket                                                                              : std_logic;                      -- width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	signal width_adapter_002_src_data                                                                                       : std_logic_vector(81 downto 0);  -- width_adapter_002:out_data -> burst_adapter_001:sink0_data
	signal width_adapter_002_src_ready                                                                                      : std_logic;                      -- burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	signal width_adapter_002_src_channel                                                                                    : std_logic_vector(14 downto 0);  -- width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	signal id_router_014_src_endofpacket                                                                                    : std_logic;                      -- id_router_014:src_endofpacket -> width_adapter_003:in_endofpacket
	signal id_router_014_src_valid                                                                                          : std_logic;                      -- id_router_014:src_valid -> width_adapter_003:in_valid
	signal id_router_014_src_startofpacket                                                                                  : std_logic;                      -- id_router_014:src_startofpacket -> width_adapter_003:in_startofpacket
	signal id_router_014_src_data                                                                                           : std_logic_vector(81 downto 0);  -- id_router_014:src_data -> width_adapter_003:in_data
	signal id_router_014_src_channel                                                                                        : std_logic_vector(14 downto 0);  -- id_router_014:src_channel -> width_adapter_003:in_channel
	signal id_router_014_src_ready                                                                                          : std_logic;                      -- width_adapter_003:in_ready -> id_router_014:src_ready
	signal width_adapter_003_src_endofpacket                                                                                : std_logic;                      -- width_adapter_003:out_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	signal width_adapter_003_src_valid                                                                                      : std_logic;                      -- width_adapter_003:out_valid -> rsp_xbar_demux_014:sink_valid
	signal width_adapter_003_src_startofpacket                                                                              : std_logic;                      -- width_adapter_003:out_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	signal width_adapter_003_src_data                                                                                       : std_logic_vector(99 downto 0);  -- width_adapter_003:out_data -> rsp_xbar_demux_014:sink_data
	signal width_adapter_003_src_ready                                                                                      : std_logic;                      -- rsp_xbar_demux_014:sink_ready -> width_adapter_003:out_ready
	signal width_adapter_003_src_channel                                                                                    : std_logic_vector(14 downto 0);  -- width_adapter_003:out_channel -> rsp_xbar_demux_014:sink_channel
	signal irq_mapper_receiver0_irq                                                                                         : std_logic;                      -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                                                         : std_logic;                      -- timer_0:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                                                         : std_logic;                      -- timer_1:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                                                                         : std_logic;                      -- de2_pio_keys4:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                                                                         : std_logic;                      -- de2_pio_toggles18:irq -> irq_mapper:receiver4_irq
	signal nios2_ht18_lemonde_streit_d_irq_irq                                                                              : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> nios2_ht18_lemonde_streit:d_irq
	signal reset_reset_n_ports_inv                                                                                          : std_logic;                      -- reset_reset_n:inv -> [rst_controller:reset_in1, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv                                     : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write:inv -> jtag_uart_0:av_write_n
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv                                      : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read:inv -> jtag_uart_0:av_read_n
	signal timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv                                                        : std_logic;                      -- timer_0_s1_translator_avalon_anti_slave_0_write:inv -> timer_0:write_n
	signal timer_1_s1_translator_avalon_anti_slave_0_write_ports_inv                                                        : std_logic;                      -- timer_1_s1_translator_avalon_anti_slave_0_write:inv -> timer_1:write_n
	signal de2_pio_toggles18_s1_translator_avalon_anti_slave_0_write_ports_inv                                              : std_logic;                      -- de2_pio_toggles18_s1_translator_avalon_anti_slave_0_write:inv -> de2_pio_toggles18:write_n
	signal de2_pio_keys4_s1_translator_avalon_anti_slave_0_write_ports_inv                                                  : std_logic;                      -- de2_pio_keys4_s1_translator_avalon_anti_slave_0_write:inv -> de2_pio_keys4:write_n
	signal de2_pio_redled18_s1_translator_avalon_anti_slave_0_write_ports_inv                                               : std_logic;                      -- de2_pio_redled18_s1_translator_avalon_anti_slave_0_write:inv -> de2_pio_redled18:write_n
	signal de2_pio_greenled9_s1_translator_avalon_anti_slave_0_write_ports_inv                                              : std_logic;                      -- de2_pio_greenled9_s1_translator_avalon_anti_slave_0_write:inv -> de2_pio_greenled9:write_n
	signal de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_write_ports_inv                                             : std_logic;                      -- de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_write:inv -> de2_pio_hex_high28:write_n
	signal de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_write_ports_inv                                              : std_logic;                      -- de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_write:inv -> de2_pio_hex_low28:write_n
	signal sdram_s1_translator_avalon_anti_slave_0_write_ports_inv                                                          : std_logic;                      -- sdram_s1_translator_avalon_anti_slave_0_write:inv -> sdram:az_wr_n
	signal sdram_s1_translator_avalon_anti_slave_0_read_ports_inv                                                           : std_logic;                      -- sdram_s1_translator_avalon_anti_slave_0_read:inv -> sdram:az_rd_n
	signal sdram_s1_translator_avalon_anti_slave_0_byteenable_ports_inv                                                     : std_logic_vector(1 downto 0);   -- sdram_s1_translator_avalon_anti_slave_0_byteenable:inv -> sdram:az_be_n
	signal rst_controller_reset_out_reset_ports_inv                                                                         : std_logic;                      -- rst_controller_reset_out_reset:inv -> [de2_pio_greenled9:reset_n, de2_pio_hex_high28:reset_n, de2_pio_hex_low28:reset_n, de2_pio_keys4:reset_n, de2_pio_redled18:reset_n, de2_pio_toggles18:reset_n, jtag_uart_0:rst_n, nios2_ht18_lemonde_streit:reset_n, p_counter:reset_n, sdram:reset_n, timer_0:reset_n, timer_1:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                                                                     : std_logic;                      -- rst_controller_001_reset_out_reset:inv -> ht18_lemonde_streit:reset_n

begin

	nios2_ht18_lemonde_streit : component nios2_ht18_lemonde_streit_nios2_ht18_lemonde_streit
		port map (
			clk                                   => up_clocks_0_sys_clk_clk,                                                                --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                                               --                   reset_n.reset_n
			d_address                             => nios2_ht18_lemonde_streit_data_master_address,                                          --               data_master.address
			d_byteenable                          => nios2_ht18_lemonde_streit_data_master_byteenable,                                       --                          .byteenable
			d_read                                => nios2_ht18_lemonde_streit_data_master_read,                                             --                          .read
			d_readdata                            => nios2_ht18_lemonde_streit_data_master_readdata,                                         --                          .readdata
			d_waitrequest                         => nios2_ht18_lemonde_streit_data_master_waitrequest,                                      --                          .waitrequest
			d_write                               => nios2_ht18_lemonde_streit_data_master_write,                                            --                          .write
			d_writedata                           => nios2_ht18_lemonde_streit_data_master_writedata,                                        --                          .writedata
			jtag_debug_module_debugaccess_to_roms => nios2_ht18_lemonde_streit_data_master_debugaccess,                                      --                          .debugaccess
			i_address                             => nios2_ht18_lemonde_streit_instruction_master_address,                                   --        instruction_master.address
			i_read                                => nios2_ht18_lemonde_streit_instruction_master_read,                                      --                          .read
			i_readdata                            => nios2_ht18_lemonde_streit_instruction_master_readdata,                                  --                          .readdata
			i_waitrequest                         => nios2_ht18_lemonde_streit_instruction_master_waitrequest,                               --                          .waitrequest
			d_irq                                 => nios2_ht18_lemonde_streit_d_irq_irq,                                                    --                     d_irq.irq
			jtag_debug_module_resetrequest        => nios2_ht18_lemonde_streit_jtag_debug_module_reset_reset,                                --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_read,        --                          .read
			jtag_debug_module_readdata            => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_write,       --                          .write
			jtag_debug_module_writedata           => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_writedata,   --                          .writedata
			no_ci_readra                          => open                                                                                    -- custom_instruction_master.readra
		);

	onchip_memory : component nios2_ht18_lemonde_streit_onchip_memory
		port map (
			clk        => up_clocks_0_sys_clk_clk,                                    --   clk1.clk
			address    => onchip_memory_s1_translator_avalon_anti_slave_0_address,    --     s1.address
			clken      => onchip_memory_s1_translator_avalon_anti_slave_0_clken,      --       .clken
			chipselect => onchip_memory_s1_translator_avalon_anti_slave_0_chipselect, --       .chipselect
			write      => onchip_memory_s1_translator_avalon_anti_slave_0_write,      --       .write
			readdata   => onchip_memory_s1_translator_avalon_anti_slave_0_readdata,   --       .readdata
			writedata  => onchip_memory_s1_translator_avalon_anti_slave_0_writedata,  --       .writedata
			byteenable => onchip_memory_s1_translator_avalon_anti_slave_0_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req                          --       .reset_req
		);

	ht18_lemonde_streit : component nios2_ht18_lemonde_streit_ht18_lemonde_streit
		port map (
			clock    => up_clocks_0_sys_clk_clk,                                                     --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,                                --         reset.reset_n
			readdata => ht18_lemonde_streit_control_slave_translator_avalon_anti_slave_0_readdata,   -- control_slave.readdata
			address  => ht18_lemonde_streit_control_slave_translator_avalon_anti_slave_0_address(0)  --              .address
		);

	jtag_uart_0 : component nios2_ht18_lemonde_streit_jtag_uart_0
		port map (
			clk            => up_clocks_0_sys_clk_clk,                                                      --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                                     --             reset.reset_n
			av_chipselect  => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address(0),      --                  .address
			av_read_n      => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			av_readdata    => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			av_write_n     => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			av_writedata   => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			av_waitrequest => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                                      --               irq.irq
		);

	timer_0 : component nios2_ht18_lemonde_streit_timer_0
		port map (
			clk        => up_clocks_0_sys_clk_clk,                                   --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                  -- reset.reset_n
			address    => timer_0_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => timer_0_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => timer_0_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => timer_0_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                                   --   irq.irq
		);

	timer_1 : component nios2_ht18_lemonde_streit_timer_1
		port map (
			clk        => up_clocks_0_sys_clk_clk,                                   --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                  -- reset.reset_n
			address    => timer_1_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => timer_1_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => timer_1_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => timer_1_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => timer_1_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver2_irq                                   --   irq.irq
		);

	p_counter : component nios2_ht18_lemonde_streit_p_counter
		port map (
			clk           => up_clocks_0_sys_clk_clk,                                              --           clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                             --         reset.reset_n
			address       => p_counter_control_slave_translator_avalon_anti_slave_0_address,       -- control_slave.address
			begintransfer => p_counter_control_slave_translator_avalon_anti_slave_0_begintransfer, --              .begintransfer
			readdata      => p_counter_control_slave_translator_avalon_anti_slave_0_readdata,      --              .readdata
			write         => p_counter_control_slave_translator_avalon_anti_slave_0_write,         --              .write
			writedata     => p_counter_control_slave_translator_avalon_anti_slave_0_writedata      --              .writedata
		);

	de2_pio_toggles18 : component nios2_ht18_lemonde_streit_de2_pio_toggles18
		port map (
			clk        => up_clocks_0_sys_clk_clk,                                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                            --               reset.reset_n
			address    => de2_pio_toggles18_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => de2_pio_toggles18_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => de2_pio_toggles18_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => de2_pio_toggles18_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => de2_pio_toggles18_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => switches18_export,                                                   -- external_connection.export
			irq        => irq_mapper_receiver4_irq                                             --                 irq.irq
		);

	de2_pio_keys4 : component nios2_ht18_lemonde_streit_de2_pio_keys4
		port map (
			clk        => up_clocks_0_sys_clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                        --               reset.reset_n
			address    => de2_pio_keys4_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => de2_pio_keys4_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => de2_pio_keys4_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => de2_pio_keys4_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => de2_pio_keys4_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => keys4_export,                                                    -- external_connection.export
			irq        => irq_mapper_receiver3_irq                                         --                 irq.irq
		);

	de2_pio_redled18 : component nios2_ht18_lemonde_streit_de2_pio_redled18
		port map (
			clk        => up_clocks_0_sys_clk_clk,                                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                           --               reset.reset_n
			address    => de2_pio_redled18_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => de2_pio_redled18_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => de2_pio_redled18_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => de2_pio_redled18_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => de2_pio_redled18_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => leds_red18_export                                                   -- external_connection.export
		);

	de2_pio_greenled9 : component nios2_ht18_lemonde_streit_de2_pio_greenled9
		port map (
			clk        => up_clocks_0_sys_clk_clk,                                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                            --               reset.reset_n
			address    => de2_pio_greenled9_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => de2_pio_greenled9_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => de2_pio_greenled9_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => de2_pio_greenled9_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => de2_pio_greenled9_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => leds_green9_export                                                   -- external_connection.export
		);

	de2_pio_hex_high28 : component nios2_ht18_lemonde_streit_de2_pio_hex_high28
		port map (
			clk        => up_clocks_0_sys_clk_clk,                                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                             --               reset.reset_n
			address    => de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => hex_high28_export                                                     -- external_connection.export
		);

	de2_pio_hex_low28 : component nios2_ht18_lemonde_streit_de2_pio_hex_high28
		port map (
			clk        => up_clocks_0_sys_clk_clk,                                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                            --               reset.reset_n
			address    => de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => hex_low28_export                                                     -- external_connection.export
		);

	sdram : component nios2_ht18_lemonde_streit_sdram
		port map (
			clk            => up_clocks_0_sys_clk_clk,                                      --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                     -- reset.reset_n
			az_addr        => sdram_s1_translator_avalon_anti_slave_0_address,              --    s1.address
			az_be_n        => sdram_s1_translator_avalon_anti_slave_0_byteenable_ports_inv, --      .byteenable_n
			az_cs          => sdram_s1_translator_avalon_anti_slave_0_chipselect,           --      .chipselect
			az_data        => sdram_s1_translator_avalon_anti_slave_0_writedata,            --      .writedata
			az_rd_n        => sdram_s1_translator_avalon_anti_slave_0_read_ports_inv,       --      .read_n
			az_wr_n        => sdram_s1_translator_avalon_anti_slave_0_write_ports_inv,      --      .write_n
			za_data        => sdram_s1_translator_avalon_anti_slave_0_readdata,             --      .readdata
			za_valid       => sdram_s1_translator_avalon_anti_slave_0_readdatavalid,        --      .readdatavalid
			za_waitrequest => sdram_s1_translator_avalon_anti_slave_0_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                              --  wire.export
			zs_ba          => sdram_wire_ba,                                                --      .export
			zs_cas_n       => sdram_wire_cas_n,                                             --      .export
			zs_cke         => sdram_wire_cke,                                               --      .export
			zs_cs_n        => sdram_wire_cs_n,                                              --      .export
			zs_dq          => sdram_wire_dq,                                                --      .export
			zs_dqm         => sdram_wire_dqm,                                               --      .export
			zs_ras_n       => sdram_wire_ras_n,                                             --      .export
			zs_we_n        => sdram_wire_we_n                                               --      .export
		);

	up_clocks_0 : component nios2_ht18_lemonde_streit_up_clocks_0
		port map (
			CLOCK_50    => clk_clk,                            --       clk_in_primary.clk
			reset       => rst_controller_002_reset_out_reset, -- clk_in_primary_reset.reset
			sys_clk     => up_clocks_0_sys_clk_clk,            --              sys_clk.clk
			sys_reset_n => open,                               --        sys_clk_reset.reset_n
			SDRAM_CLK   => sdram_clk_clk                       --            sdram_clk.clk
		);

	sram : component nios2_ht18_lemonde_streit_sram
		port map (
			clk           => up_clocks_0_sys_clk_clk,                                             --        clock_reset.clk
			reset         => rst_controller_reset_out_reset,                                      --  clock_reset_reset.reset
			SRAM_DQ       => sram_wire_DQ,                                                        -- external_interface.export
			SRAM_ADDR     => sram_wire_ADDR,                                                      --                   .export
			SRAM_LB_N     => sram_wire_LB_N,                                                      --                   .export
			SRAM_UB_N     => sram_wire_UB_N,                                                      --                   .export
			SRAM_CE_N     => sram_wire_CE_N,                                                      --                   .export
			SRAM_OE_N     => sram_wire_OE_N,                                                      --                   .export
			SRAM_WE_N     => sram_wire_WE_N,                                                      --                   .export
			address       => sram_avalon_sram_slave_translator_avalon_anti_slave_0_address,       --  avalon_sram_slave.address
			byteenable    => sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable,    --                   .byteenable
			read          => sram_avalon_sram_slave_translator_avalon_anti_slave_0_read,          --                   .read
			write         => sram_avalon_sram_slave_translator_avalon_anti_slave_0_write,         --                   .write
			writedata     => sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata,     --                   .writedata
			readdata      => sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata,      --                   .readdata
			readdatavalid => sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid  --                   .readdatavalid
		);

	nios2_ht18_lemonde_streit_data_master_translator : component nios2_ht18_lemonde_streit_nios2_ht18_lemonde_streit_data_master_translator
		generic map (
			AV_ADDRESS_W                => 25,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 25,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 1
		)
		port map (
			clk                      => up_clocks_0_sys_clk_clk,                                                                  --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                                           --                     reset.reset
			uav_address              => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => nios2_ht18_lemonde_streit_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => nios2_ht18_lemonde_streit_data_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => nios2_ht18_lemonde_streit_data_master_byteenable,                                         --                          .byteenable
			av_read                  => nios2_ht18_lemonde_streit_data_master_read,                                               --                          .read
			av_readdata              => nios2_ht18_lemonde_streit_data_master_readdata,                                           --                          .readdata
			av_write                 => nios2_ht18_lemonde_streit_data_master_write,                                              --                          .write
			av_writedata             => nios2_ht18_lemonde_streit_data_master_writedata,                                          --                          .writedata
			av_debugaccess           => nios2_ht18_lemonde_streit_data_master_debugaccess,                                        --                          .debugaccess
			av_burstcount            => "1",                                                                                      --               (terminated)
			av_beginbursttransfer    => '0',                                                                                      --               (terminated)
			av_begintransfer         => '0',                                                                                      --               (terminated)
			av_chipselect            => '0',                                                                                      --               (terminated)
			av_readdatavalid         => open,                                                                                     --               (terminated)
			av_lock                  => '0',                                                                                      --               (terminated)
			uav_clken                => open,                                                                                     --               (terminated)
			av_clken                 => '1',                                                                                      --               (terminated)
			uav_response             => "00",                                                                                     --               (terminated)
			av_response              => open,                                                                                     --               (terminated)
			uav_writeresponserequest => open,                                                                                     --               (terminated)
			uav_writeresponsevalid   => '0',                                                                                      --               (terminated)
			av_writeresponserequest  => '0',                                                                                      --               (terminated)
			av_writeresponsevalid    => open                                                                                      --               (terminated)
		);

	nios2_ht18_lemonde_streit_instruction_master_translator : component nios2_ht18_lemonde_streit_nios2_ht18_lemonde_streit_instruction_master_translator
		generic map (
			AV_ADDRESS_W                => 25,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 25,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 1,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => up_clocks_0_sys_clk_clk,                                                                         --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                                                  --                     reset.reset
			uav_address              => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => nios2_ht18_lemonde_streit_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => nios2_ht18_lemonde_streit_instruction_master_waitrequest,                                        --                          .waitrequest
			av_read                  => nios2_ht18_lemonde_streit_instruction_master_read,                                               --                          .read
			av_readdata              => nios2_ht18_lemonde_streit_instruction_master_readdata,                                           --                          .readdata
			av_burstcount            => "1",                                                                                             --               (terminated)
			av_byteenable            => "1111",                                                                                          --               (terminated)
			av_beginbursttransfer    => '0',                                                                                             --               (terminated)
			av_begintransfer         => '0',                                                                                             --               (terminated)
			av_chipselect            => '0',                                                                                             --               (terminated)
			av_readdatavalid         => open,                                                                                            --               (terminated)
			av_write                 => '0',                                                                                             --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                                              --               (terminated)
			av_lock                  => '0',                                                                                             --               (terminated)
			av_debugaccess           => '0',                                                                                             --               (terminated)
			uav_clken                => open,                                                                                            --               (terminated)
			av_clken                 => '1',                                                                                             --               (terminated)
			uav_response             => "00",                                                                                            --               (terminated)
			av_response              => open,                                                                                            --               (terminated)
			uav_writeresponserequest => open,                                                                                            --               (terminated)
			uav_writeresponsevalid   => '0',                                                                                             --               (terminated)
			av_writeresponserequest  => '0',                                                                                             --               (terminated)
			av_writeresponsevalid    => open                                                                                             --               (terminated)
		);

	onchip_memory_s1_translator : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator
		generic map (
			AV_ADDRESS_W                   => 13,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => up_clocks_0_sys_clk_clk,                                                     --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                              --                    reset.reset
			uav_address              => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => onchip_memory_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => onchip_memory_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => onchip_memory_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => onchip_memory_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => onchip_memory_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect            => onchip_memory_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_clken                 => onchip_memory_s1_translator_avalon_anti_slave_0_clken,                       --                         .clken
			av_read                  => open,                                                                        --              (terminated)
			av_begintransfer         => open,                                                                        --              (terminated)
			av_beginbursttransfer    => open,                                                                        --              (terminated)
			av_burstcount            => open,                                                                        --              (terminated)
			av_readdatavalid         => '0',                                                                         --              (terminated)
			av_waitrequest           => '0',                                                                         --              (terminated)
			av_writebyteenable       => open,                                                                        --              (terminated)
			av_lock                  => open,                                                                        --              (terminated)
			uav_clken                => '0',                                                                         --              (terminated)
			av_debugaccess           => open,                                                                        --              (terminated)
			av_outputenable          => open,                                                                        --              (terminated)
			uav_response             => open,                                                                        --              (terminated)
			av_response              => "00",                                                                        --              (terminated)
			uav_writeresponserequest => '0',                                                                         --              (terminated)
			uav_writeresponsevalid   => open,                                                                        --              (terminated)
			av_writeresponserequest  => open,                                                                        --              (terminated)
			av_writeresponsevalid    => '0'                                                                          --              (terminated)
		);

	ht18_lemonde_streit_control_slave_translator : component nios2_ht18_lemonde_streit_ht18_lemonde_streit_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => up_clocks_0_sys_clk_clk,                                                                      --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                           --                    reset.reset
			uav_address              => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => ht18_lemonde_streit_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => ht18_lemonde_streit_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                                         --              (terminated)
			av_read                  => open,                                                                                         --              (terminated)
			av_writedata             => open,                                                                                         --              (terminated)
			av_begintransfer         => open,                                                                                         --              (terminated)
			av_beginbursttransfer    => open,                                                                                         --              (terminated)
			av_burstcount            => open,                                                                                         --              (terminated)
			av_byteenable            => open,                                                                                         --              (terminated)
			av_readdatavalid         => '0',                                                                                          --              (terminated)
			av_waitrequest           => '0',                                                                                          --              (terminated)
			av_writebyteenable       => open,                                                                                         --              (terminated)
			av_lock                  => open,                                                                                         --              (terminated)
			av_chipselect            => open,                                                                                         --              (terminated)
			av_clken                 => open,                                                                                         --              (terminated)
			uav_clken                => '0',                                                                                          --              (terminated)
			av_debugaccess           => open,                                                                                         --              (terminated)
			av_outputenable          => open,                                                                                         --              (terminated)
			uav_response             => open,                                                                                         --              (terminated)
			av_response              => "00",                                                                                         --              (terminated)
			uav_writeresponserequest => '0',                                                                                          --              (terminated)
			uav_writeresponsevalid   => open,                                                                                         --              (terminated)
			av_writeresponserequest  => open,                                                                                         --              (terminated)
			av_writeresponsevalid    => '0'                                                                                           --              (terminated)
		);

	jtag_uart_0_avalon_jtag_slave_translator : component nios2_ht18_lemonde_streit_jtag_uart_0_avalon_jtag_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => up_clocks_0_sys_clk_clk,                                                                  --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                           --                    reset.reset
			uav_address              => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest           => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                                     --              (terminated)
			av_burstcount            => open,                                                                                     --              (terminated)
			av_byteenable            => open,                                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                                     --              (terminated)
			av_lock                  => open,                                                                                     --              (terminated)
			av_clken                 => open,                                                                                     --              (terminated)
			uav_clken                => '0',                                                                                      --              (terminated)
			av_debugaccess           => open,                                                                                     --              (terminated)
			av_outputenable          => open,                                                                                     --              (terminated)
			uav_response             => open,                                                                                     --              (terminated)
			av_response              => "00",                                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                                       --              (terminated)
		);

	nios2_ht18_lemonde_streit_jtag_debug_module_translator : component nios2_ht18_lemonde_streit_nios2_ht18_lemonde_streit_jtag_debug_module_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => up_clocks_0_sys_clk_clk,                                                                                --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                                         --                    reset.reset
			uav_address              => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                                                   --              (terminated)
			av_burstcount            => open,                                                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                                                   --              (terminated)
			av_lock                  => open,                                                                                                   --              (terminated)
			av_chipselect            => open,                                                                                                   --              (terminated)
			av_clken                 => open,                                                                                                   --              (terminated)
			uav_clken                => '0',                                                                                                    --              (terminated)
			av_outputenable          => open,                                                                                                   --              (terminated)
			uav_response             => open,                                                                                                   --              (terminated)
			av_response              => "00",                                                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                                                     --              (terminated)
		);

	timer_0_s1_translator : component nios2_ht18_lemonde_streit_timer_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => up_clocks_0_sys_clk_clk,                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => timer_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => timer_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => timer_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => timer_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => timer_0_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	timer_1_s1_translator : component nios2_ht18_lemonde_streit_timer_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => up_clocks_0_sys_clk_clk,                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => timer_1_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => timer_1_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => timer_1_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => timer_1_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => timer_1_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	p_counter_control_slave_translator : component nios2_ht18_lemonde_streit_p_counter_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 5,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => up_clocks_0_sys_clk_clk,                                                            --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                     --                    reset.reset
			uav_address              => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => p_counter_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => p_counter_control_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => p_counter_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => p_counter_control_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer         => p_counter_control_slave_translator_avalon_anti_slave_0_begintransfer,               --                         .begintransfer
			av_read                  => open,                                                                               --              (terminated)
			av_beginbursttransfer    => open,                                                                               --              (terminated)
			av_burstcount            => open,                                                                               --              (terminated)
			av_byteenable            => open,                                                                               --              (terminated)
			av_readdatavalid         => '0',                                                                                --              (terminated)
			av_waitrequest           => '0',                                                                                --              (terminated)
			av_writebyteenable       => open,                                                                               --              (terminated)
			av_lock                  => open,                                                                               --              (terminated)
			av_chipselect            => open,                                                                               --              (terminated)
			av_clken                 => open,                                                                               --              (terminated)
			uav_clken                => '0',                                                                                --              (terminated)
			av_debugaccess           => open,                                                                               --              (terminated)
			av_outputenable          => open,                                                                               --              (terminated)
			uav_response             => open,                                                                               --              (terminated)
			av_response              => "00",                                                                               --              (terminated)
			uav_writeresponserequest => '0',                                                                                --              (terminated)
			uav_writeresponsevalid   => open,                                                                               --              (terminated)
			av_writeresponserequest  => open,                                                                               --              (terminated)
			av_writeresponsevalid    => '0'                                                                                 --              (terminated)
		);

	de2_pio_toggles18_s1_translator : component nios2_ht18_lemonde_streit_de2_pio_toggles18_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => up_clocks_0_sys_clk_clk,                                                         --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                  --                    reset.reset
			uav_address              => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => de2_pio_toggles18_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => de2_pio_toggles18_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => de2_pio_toggles18_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => de2_pio_toggles18_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => de2_pio_toggles18_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                            --              (terminated)
			av_begintransfer         => open,                                                                            --              (terminated)
			av_beginbursttransfer    => open,                                                                            --              (terminated)
			av_burstcount            => open,                                                                            --              (terminated)
			av_byteenable            => open,                                                                            --              (terminated)
			av_readdatavalid         => '0',                                                                             --              (terminated)
			av_waitrequest           => '0',                                                                             --              (terminated)
			av_writebyteenable       => open,                                                                            --              (terminated)
			av_lock                  => open,                                                                            --              (terminated)
			av_clken                 => open,                                                                            --              (terminated)
			uav_clken                => '0',                                                                             --              (terminated)
			av_debugaccess           => open,                                                                            --              (terminated)
			av_outputenable          => open,                                                                            --              (terminated)
			uav_response             => open,                                                                            --              (terminated)
			av_response              => "00",                                                                            --              (terminated)
			uav_writeresponserequest => '0',                                                                             --              (terminated)
			uav_writeresponsevalid   => open,                                                                            --              (terminated)
			av_writeresponserequest  => open,                                                                            --              (terminated)
			av_writeresponsevalid    => '0'                                                                              --              (terminated)
		);

	de2_pio_keys4_s1_translator : component nios2_ht18_lemonde_streit_de2_pio_toggles18_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => up_clocks_0_sys_clk_clk,                                                     --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                              --                    reset.reset
			uav_address              => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => de2_pio_keys4_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => de2_pio_keys4_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => de2_pio_keys4_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => de2_pio_keys4_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => de2_pio_keys4_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                        --              (terminated)
			av_begintransfer         => open,                                                                        --              (terminated)
			av_beginbursttransfer    => open,                                                                        --              (terminated)
			av_burstcount            => open,                                                                        --              (terminated)
			av_byteenable            => open,                                                                        --              (terminated)
			av_readdatavalid         => '0',                                                                         --              (terminated)
			av_waitrequest           => '0',                                                                         --              (terminated)
			av_writebyteenable       => open,                                                                        --              (terminated)
			av_lock                  => open,                                                                        --              (terminated)
			av_clken                 => open,                                                                        --              (terminated)
			uav_clken                => '0',                                                                         --              (terminated)
			av_debugaccess           => open,                                                                        --              (terminated)
			av_outputenable          => open,                                                                        --              (terminated)
			uav_response             => open,                                                                        --              (terminated)
			av_response              => "00",                                                                        --              (terminated)
			uav_writeresponserequest => '0',                                                                         --              (terminated)
			uav_writeresponsevalid   => open,                                                                        --              (terminated)
			av_writeresponserequest  => open,                                                                        --              (terminated)
			av_writeresponsevalid    => '0'                                                                          --              (terminated)
		);

	de2_pio_redled18_s1_translator : component nios2_ht18_lemonde_streit_de2_pio_toggles18_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => up_clocks_0_sys_clk_clk,                                                        --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                 --                    reset.reset
			uav_address              => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => de2_pio_redled18_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => de2_pio_redled18_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => de2_pio_redled18_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => de2_pio_redled18_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => de2_pio_redled18_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                           --              (terminated)
			av_begintransfer         => open,                                                                           --              (terminated)
			av_beginbursttransfer    => open,                                                                           --              (terminated)
			av_burstcount            => open,                                                                           --              (terminated)
			av_byteenable            => open,                                                                           --              (terminated)
			av_readdatavalid         => '0',                                                                            --              (terminated)
			av_waitrequest           => '0',                                                                            --              (terminated)
			av_writebyteenable       => open,                                                                           --              (terminated)
			av_lock                  => open,                                                                           --              (terminated)
			av_clken                 => open,                                                                           --              (terminated)
			uav_clken                => '0',                                                                            --              (terminated)
			av_debugaccess           => open,                                                                           --              (terminated)
			av_outputenable          => open,                                                                           --              (terminated)
			uav_response             => open,                                                                           --              (terminated)
			av_response              => "00",                                                                           --              (terminated)
			uav_writeresponserequest => '0',                                                                            --              (terminated)
			uav_writeresponsevalid   => open,                                                                           --              (terminated)
			av_writeresponserequest  => open,                                                                           --              (terminated)
			av_writeresponsevalid    => '0'                                                                             --              (terminated)
		);

	de2_pio_greenled9_s1_translator : component nios2_ht18_lemonde_streit_de2_pio_toggles18_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => up_clocks_0_sys_clk_clk,                                                         --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                  --                    reset.reset
			uav_address              => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => de2_pio_greenled9_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => de2_pio_greenled9_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => de2_pio_greenled9_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => de2_pio_greenled9_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => de2_pio_greenled9_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                            --              (terminated)
			av_begintransfer         => open,                                                                            --              (terminated)
			av_beginbursttransfer    => open,                                                                            --              (terminated)
			av_burstcount            => open,                                                                            --              (terminated)
			av_byteenable            => open,                                                                            --              (terminated)
			av_readdatavalid         => '0',                                                                             --              (terminated)
			av_waitrequest           => '0',                                                                             --              (terminated)
			av_writebyteenable       => open,                                                                            --              (terminated)
			av_lock                  => open,                                                                            --              (terminated)
			av_clken                 => open,                                                                            --              (terminated)
			uav_clken                => '0',                                                                             --              (terminated)
			av_debugaccess           => open,                                                                            --              (terminated)
			av_outputenable          => open,                                                                            --              (terminated)
			uav_response             => open,                                                                            --              (terminated)
			av_response              => "00",                                                                            --              (terminated)
			uav_writeresponserequest => '0',                                                                             --              (terminated)
			uav_writeresponsevalid   => open,                                                                            --              (terminated)
			av_writeresponserequest  => open,                                                                            --              (terminated)
			av_writeresponsevalid    => '0'                                                                              --              (terminated)
		);

	de2_pio_hex_high28_s1_translator : component nios2_ht18_lemonde_streit_de2_pio_toggles18_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => up_clocks_0_sys_clk_clk,                                                          --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                   --                    reset.reset
			uav_address              => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                             --              (terminated)
			av_begintransfer         => open,                                                                             --              (terminated)
			av_beginbursttransfer    => open,                                                                             --              (terminated)
			av_burstcount            => open,                                                                             --              (terminated)
			av_byteenable            => open,                                                                             --              (terminated)
			av_readdatavalid         => '0',                                                                              --              (terminated)
			av_waitrequest           => '0',                                                                              --              (terminated)
			av_writebyteenable       => open,                                                                             --              (terminated)
			av_lock                  => open,                                                                             --              (terminated)
			av_clken                 => open,                                                                             --              (terminated)
			uav_clken                => '0',                                                                              --              (terminated)
			av_debugaccess           => open,                                                                             --              (terminated)
			av_outputenable          => open,                                                                             --              (terminated)
			uav_response             => open,                                                                             --              (terminated)
			av_response              => "00",                                                                             --              (terminated)
			uav_writeresponserequest => '0',                                                                              --              (terminated)
			uav_writeresponsevalid   => open,                                                                             --              (terminated)
			av_writeresponserequest  => open,                                                                             --              (terminated)
			av_writeresponsevalid    => '0'                                                                               --              (terminated)
		);

	de2_pio_hex_low28_s1_translator : component nios2_ht18_lemonde_streit_de2_pio_toggles18_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => up_clocks_0_sys_clk_clk,                                                         --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                  --                    reset.reset
			uav_address              => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                            --              (terminated)
			av_begintransfer         => open,                                                                            --              (terminated)
			av_beginbursttransfer    => open,                                                                            --              (terminated)
			av_burstcount            => open,                                                                            --              (terminated)
			av_byteenable            => open,                                                                            --              (terminated)
			av_readdatavalid         => '0',                                                                             --              (terminated)
			av_waitrequest           => '0',                                                                             --              (terminated)
			av_writebyteenable       => open,                                                                            --              (terminated)
			av_lock                  => open,                                                                            --              (terminated)
			av_clken                 => open,                                                                            --              (terminated)
			uav_clken                => '0',                                                                             --              (terminated)
			av_debugaccess           => open,                                                                            --              (terminated)
			av_outputenable          => open,                                                                            --              (terminated)
			uav_response             => open,                                                                            --              (terminated)
			av_response              => "00",                                                                            --              (terminated)
			uav_writeresponserequest => '0',                                                                             --              (terminated)
			uav_writeresponsevalid   => open,                                                                            --              (terminated)
			av_writeresponserequest  => open,                                                                            --              (terminated)
			av_writeresponsevalid    => '0'                                                                              --              (terminated)
		);

	sram_avalon_sram_slave_translator : component nios2_ht18_lemonde_streit_sram_avalon_sram_slave_translator
		generic map (
			AV_ADDRESS_W                   => 18,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => up_clocks_0_sys_clk_clk,                                                           --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                    --                    reset.reset
			uav_address              => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sram_avalon_sram_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sram_avalon_sram_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => sram_avalon_sram_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_begintransfer         => open,                                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                                              --              (terminated)
			av_burstcount            => open,                                                                              --              (terminated)
			av_waitrequest           => '0',                                                                               --              (terminated)
			av_writebyteenable       => open,                                                                              --              (terminated)
			av_lock                  => open,                                                                              --              (terminated)
			av_chipselect            => open,                                                                              --              (terminated)
			av_clken                 => open,                                                                              --              (terminated)
			uav_clken                => '0',                                                                               --              (terminated)
			av_debugaccess           => open,                                                                              --              (terminated)
			av_outputenable          => open,                                                                              --              (terminated)
			uav_response             => open,                                                                              --              (terminated)
			av_response              => "00",                                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                                              --              (terminated)
			av_writeresponserequest  => open,                                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                                --              (terminated)
		);

	sdram_s1_translator : component nios2_ht18_lemonde_streit_sdram_s1_translator
		generic map (
			AV_ADDRESS_W                   => 22,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => up_clocks_0_sys_clk_clk,                                             --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                      --                    reset.reset
			uav_address              => sdram_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sdram_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sdram_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sdram_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sdram_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => sdram_s1_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => sdram_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sdram_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => sdram_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => sdram_s1_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => sdram_s1_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => sdram_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                --              (terminated)
			av_beginbursttransfer    => open,                                                                --              (terminated)
			av_burstcount            => open,                                                                --              (terminated)
			av_writebyteenable       => open,                                                                --              (terminated)
			av_lock                  => open,                                                                --              (terminated)
			av_clken                 => open,                                                                --              (terminated)
			uav_clken                => '0',                                                                 --              (terminated)
			av_debugaccess           => open,                                                                --              (terminated)
			av_outputenable          => open,                                                                --              (terminated)
			uav_response             => open,                                                                --              (terminated)
			av_response              => "00",                                                                --              (terminated)
			uav_writeresponserequest => '0',                                                                 --              (terminated)
			uav_writeresponsevalid   => open,                                                                --              (terminated)
			av_writeresponserequest  => open,                                                                --              (terminated)
			av_writeresponsevalid    => '0'                                                                  --              (terminated)
		);

	nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_BEGIN_BURST           => 80,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			PKT_BURST_TYPE_H          => 77,
			PKT_BURST_TYPE_L          => 76,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_TRANS_EXCLUSIVE       => 66,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_THREAD_ID_H           => 90,
			PKT_THREAD_ID_L           => 90,
			PKT_CACHE_H               => 97,
			PKT_CACHE_L               => 94,
			PKT_DATA_SIDEBAND_H       => 79,
			PKT_DATA_SIDEBAND_L       => 79,
			PKT_QOS_H                 => 81,
			PKT_QOS_L                 => 81,
			PKT_ADDR_SIDEBAND_H       => 78,
			PKT_ADDR_SIDEBAND_L       => 78,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			ST_DATA_W                 => 100,
			ST_CHANNEL_W              => 15,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                           --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                    -- clk_reset.reset
			av_address              => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_src_valid,                                                                            --        rp.valid
			rp_data                 => rsp_xbar_mux_src_data,                                                                             --          .data
			rp_channel              => rsp_xbar_mux_src_channel,                                                                          --          .channel
			rp_startofpacket        => rsp_xbar_mux_src_startofpacket,                                                                    --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_src_endofpacket,                                                                      --          .endofpacket
			rp_ready                => rsp_xbar_mux_src_ready,                                                                            --          .ready
			av_response             => open,                                                                                              -- (terminated)
			av_writeresponserequest => '0',                                                                                               -- (terminated)
			av_writeresponsevalid   => open                                                                                               -- (terminated)
		);

	nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_BEGIN_BURST           => 80,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			PKT_BURST_TYPE_H          => 77,
			PKT_BURST_TYPE_L          => 76,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_TRANS_EXCLUSIVE       => 66,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_THREAD_ID_H           => 90,
			PKT_THREAD_ID_L           => 90,
			PKT_CACHE_H               => 97,
			PKT_CACHE_L               => 94,
			PKT_DATA_SIDEBAND_H       => 79,
			PKT_DATA_SIDEBAND_L       => 79,
			PKT_QOS_H                 => 81,
			PKT_QOS_L                 => 81,
			PKT_ADDR_SIDEBAND_H       => 78,
			PKT_ADDR_SIDEBAND_L       => 78,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			ST_DATA_W                 => 100,
			ST_CHANNEL_W              => 15,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 1,
			BURSTWRAP_VALUE           => 3,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                                  --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                           -- clk_reset.reset
			av_address              => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_001_src_valid,                                                                               --        rp.valid
			rp_data                 => rsp_xbar_mux_001_src_data,                                                                                --          .data
			rp_channel              => rsp_xbar_mux_001_src_channel,                                                                             --          .channel
			rp_startofpacket        => rsp_xbar_mux_001_src_startofpacket,                                                                       --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_001_src_endofpacket,                                                                         --          .endofpacket
			rp_ready                => rsp_xbar_mux_001_src_ready,                                                                               --          .ready
			av_response             => open,                                                                                                     -- (terminated)
			av_writeresponserequest => '0',                                                                                                      -- (terminated)
			av_writeresponsevalid   => open                                                                                                      -- (terminated)
		);

	onchip_memory_s1_translator_avalon_universal_slave_0_agent : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 15,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                               --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                        --       clk_reset.reset
			m0_address              => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_src_ready,                                                                --              cp.ready
			cp_valid                => cmd_xbar_mux_src_valid,                                                                --                .valid
			cp_data                 => cmd_xbar_mux_src_data,                                                                 --                .data
			cp_startofpacket        => cmd_xbar_mux_src_startofpacket,                                                        --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_src_endofpacket,                                                          --                .endofpacket
			cp_channel              => cmd_xbar_mux_src_channel,                                                              --                .channel
			rf_sink_ready           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                  --     (terminated)
			m0_writeresponserequest => open,                                                                                  --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                    --     (terminated)
		);

	onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                               --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			in_data           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                  -- (terminated)
			csr_read          => '0',                                                                                   -- (terminated)
			csr_write         => '0',                                                                                   -- (terminated)
			csr_readdata      => open,                                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                    -- (terminated)
			almost_full_data  => open,                                                                                  -- (terminated)
			almost_empty_data => open,                                                                                  -- (terminated)
			in_empty          => '0',                                                                                   -- (terminated)
			out_empty         => open,                                                                                  -- (terminated)
			in_error          => '0',                                                                                   -- (terminated)
			out_error         => open,                                                                                  -- (terminated)
			in_channel        => '0',                                                                                   -- (terminated)
			out_channel       => open                                                                                   -- (terminated)
		);

	ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 15,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                                --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                                     --       clk_reset.reset
			m0_address              => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_src1_ready,                                                                              --              cp.ready
			cp_valid                => cmd_xbar_demux_src1_valid,                                                                              --                .valid
			cp_data                 => cmd_xbar_demux_src1_data,                                                                               --                .data
			cp_startofpacket        => cmd_xbar_demux_src1_startofpacket,                                                                      --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_src1_endofpacket,                                                                        --                .endofpacket
			cp_channel              => cmd_xbar_demux_src1_channel,                                                                            --                .channel
			rf_sink_ready           => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                   --     (terminated)
			m0_writeresponserequest => open,                                                                                                   --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                     --     (terminated)
		);

	ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                                --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                                     -- clk_reset.reset
			in_data           => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                   -- (terminated)
			csr_read          => '0',                                                                                                    -- (terminated)
			csr_write         => '0',                                                                                                    -- (terminated)
			csr_readdata      => open,                                                                                                   -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                     -- (terminated)
			almost_full_data  => open,                                                                                                   -- (terminated)
			almost_empty_data => open,                                                                                                   -- (terminated)
			in_empty          => '0',                                                                                                    -- (terminated)
			out_empty         => open,                                                                                                   -- (terminated)
			in_error          => '0',                                                                                                    -- (terminated)
			out_error         => open,                                                                                                   -- (terminated)
			in_channel        => '0',                                                                                                    -- (terminated)
			out_channel       => open                                                                                                    -- (terminated)
		);

	jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 15,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                     --       clk_reset.reset
			m0_address              => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_src2_ready,                                                                          --              cp.ready
			cp_valid                => cmd_xbar_demux_src2_valid,                                                                          --                .valid
			cp_data                 => cmd_xbar_demux_src2_data,                                                                           --                .data
			cp_startofpacket        => cmd_xbar_demux_src2_startofpacket,                                                                  --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_src2_endofpacket,                                                                    --                .endofpacket
			cp_channel              => cmd_xbar_demux_src2_channel,                                                                        --                .channel
			rf_sink_ready           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                 --     (terminated)
		);

	jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                     -- clk_reset.reset
			in_data           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                               -- (terminated)
			csr_read          => '0',                                                                                                -- (terminated)
			csr_write         => '0',                                                                                                -- (terminated)
			csr_readdata      => open,                                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                 -- (terminated)
			almost_full_data  => open,                                                                                               -- (terminated)
			almost_empty_data => open,                                                                                               -- (terminated)
			in_empty          => '0',                                                                                                -- (terminated)
			out_empty         => open,                                                                                               -- (terminated)
			in_error          => '0',                                                                                                -- (terminated)
			out_error         => open,                                                                                               -- (terminated)
			in_channel        => '0',                                                                                                -- (terminated)
			out_channel       => open                                                                                                -- (terminated)
		);

	nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 15,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                                          --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                                   --       clk_reset.reset
			m0_address              => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_003_src_ready,                                                                                       --              cp.ready
			cp_valid                => cmd_xbar_mux_003_src_valid,                                                                                       --                .valid
			cp_data                 => cmd_xbar_mux_003_src_data,                                                                                        --                .data
			cp_startofpacket        => cmd_xbar_mux_003_src_startofpacket,                                                                               --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_003_src_endofpacket,                                                                                 --                .endofpacket
			cp_channel              => cmd_xbar_mux_003_src_channel,                                                                                     --                .channel
			rf_sink_ready           => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                               --     (terminated)
		);

	nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                                          --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                                   -- clk_reset.reset
			in_data           => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                             -- (terminated)
			csr_read          => '0',                                                                                                              -- (terminated)
			csr_write         => '0',                                                                                                              -- (terminated)
			csr_readdata      => open,                                                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                               -- (terminated)
			almost_full_data  => open,                                                                                                             -- (terminated)
			almost_empty_data => open,                                                                                                             -- (terminated)
			in_empty          => '0',                                                                                                              -- (terminated)
			out_empty         => open,                                                                                                             -- (terminated)
			in_error          => '0',                                                                                                              -- (terminated)
			out_error         => open,                                                                                                             -- (terminated)
			in_channel        => '0',                                                                                                              -- (terminated)
			out_channel       => open                                                                                                              -- (terminated)
		);

	timer_0_s1_translator_avalon_universal_slave_0_agent : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 15,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_src4_ready,                                                       --              cp.ready
			cp_valid                => cmd_xbar_demux_src4_valid,                                                       --                .valid
			cp_data                 => cmd_xbar_demux_src4_data,                                                        --                .data
			cp_startofpacket        => cmd_xbar_demux_src4_startofpacket,                                               --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_src4_endofpacket,                                                 --                .endofpacket
			cp_channel              => cmd_xbar_demux_src4_channel,                                                     --                .channel
			rf_sink_ready           => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	timer_1_s1_translator_avalon_universal_slave_0_agent : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 15,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_src5_ready,                                                       --              cp.ready
			cp_valid                => cmd_xbar_demux_src5_valid,                                                       --                .valid
			cp_data                 => cmd_xbar_demux_src5_data,                                                        --                .data
			cp_startofpacket        => cmd_xbar_demux_src5_startofpacket,                                               --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_src5_endofpacket,                                                 --                .endofpacket
			cp_channel              => cmd_xbar_demux_src5_channel,                                                     --                .channel
			rf_sink_ready           => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	p_counter_control_slave_translator_avalon_universal_slave_0_agent : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 15,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                      --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                               --       clk_reset.reset
			m0_address              => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => p_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_src6_ready,                                                                    --              cp.ready
			cp_valid                => cmd_xbar_demux_src6_valid,                                                                    --                .valid
			cp_data                 => cmd_xbar_demux_src6_data,                                                                     --                .data
			cp_startofpacket        => cmd_xbar_demux_src6_startofpacket,                                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_src6_endofpacket,                                                              --                .endofpacket
			cp_channel              => cmd_xbar_demux_src6_channel,                                                                  --                .channel
			rf_sink_ready           => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                         --     (terminated)
			m0_writeresponserequest => open,                                                                                         --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                           --     (terminated)
		);

	p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                      --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                               -- clk_reset.reset
			in_data           => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                         -- (terminated)
			csr_read          => '0',                                                                                          -- (terminated)
			csr_write         => '0',                                                                                          -- (terminated)
			csr_readdata      => open,                                                                                         -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                           -- (terminated)
			almost_full_data  => open,                                                                                         -- (terminated)
			almost_empty_data => open,                                                                                         -- (terminated)
			in_empty          => '0',                                                                                          -- (terminated)
			out_empty         => open,                                                                                         -- (terminated)
			in_error          => '0',                                                                                          -- (terminated)
			out_error         => open,                                                                                         -- (terminated)
			in_channel        => '0',                                                                                          -- (terminated)
			out_channel       => open                                                                                          -- (terminated)
		);

	de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 15,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                   --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                            --       clk_reset.reset
			m0_address              => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_src7_ready,                                                                 --              cp.ready
			cp_valid                => cmd_xbar_demux_src7_valid,                                                                 --                .valid
			cp_data                 => cmd_xbar_demux_src7_data,                                                                  --                .data
			cp_startofpacket        => cmd_xbar_demux_src7_startofpacket,                                                         --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_src7_endofpacket,                                                           --                .endofpacket
			cp_channel              => cmd_xbar_demux_src7_channel,                                                               --                .channel
			rf_sink_ready           => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                      --     (terminated)
			m0_writeresponserequest => open,                                                                                      --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                        --     (terminated)
		);

	de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                   --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			in_data           => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                      -- (terminated)
			csr_read          => '0',                                                                                       -- (terminated)
			csr_write         => '0',                                                                                       -- (terminated)
			csr_readdata      => open,                                                                                      -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                        -- (terminated)
			almost_full_data  => open,                                                                                      -- (terminated)
			almost_empty_data => open,                                                                                      -- (terminated)
			in_empty          => '0',                                                                                       -- (terminated)
			out_empty         => open,                                                                                      -- (terminated)
			in_error          => '0',                                                                                       -- (terminated)
			out_error         => open,                                                                                      -- (terminated)
			in_channel        => '0',                                                                                       -- (terminated)
			out_channel       => open                                                                                       -- (terminated)
		);

	de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 15,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                               --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                        --       clk_reset.reset
			m0_address              => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_src8_ready,                                                             --              cp.ready
			cp_valid                => cmd_xbar_demux_src8_valid,                                                             --                .valid
			cp_data                 => cmd_xbar_demux_src8_data,                                                              --                .data
			cp_startofpacket        => cmd_xbar_demux_src8_startofpacket,                                                     --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_src8_endofpacket,                                                       --                .endofpacket
			cp_channel              => cmd_xbar_demux_src8_channel,                                                           --                .channel
			rf_sink_ready           => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                  --     (terminated)
			m0_writeresponserequest => open,                                                                                  --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                    --     (terminated)
		);

	de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                               --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			in_data           => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                  -- (terminated)
			csr_read          => '0',                                                                                   -- (terminated)
			csr_write         => '0',                                                                                   -- (terminated)
			csr_readdata      => open,                                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                    -- (terminated)
			almost_full_data  => open,                                                                                  -- (terminated)
			almost_empty_data => open,                                                                                  -- (terminated)
			in_empty          => '0',                                                                                   -- (terminated)
			out_empty         => open,                                                                                  -- (terminated)
			in_error          => '0',                                                                                   -- (terminated)
			out_error         => open,                                                                                  -- (terminated)
			in_channel        => '0',                                                                                   -- (terminated)
			out_channel       => open                                                                                   -- (terminated)
		);

	de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 15,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                  --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                           --       clk_reset.reset
			m0_address              => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_src9_ready,                                                                --              cp.ready
			cp_valid                => cmd_xbar_demux_src9_valid,                                                                --                .valid
			cp_data                 => cmd_xbar_demux_src9_data,                                                                 --                .data
			cp_startofpacket        => cmd_xbar_demux_src9_startofpacket,                                                        --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_src9_endofpacket,                                                          --                .endofpacket
			cp_channel              => cmd_xbar_demux_src9_channel,                                                              --                .channel
			rf_sink_ready           => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                     --     (terminated)
			m0_writeresponserequest => open,                                                                                     --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                       --     (terminated)
		);

	de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                  --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                           -- clk_reset.reset
			in_data           => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                     -- (terminated)
			csr_read          => '0',                                                                                      -- (terminated)
			csr_write         => '0',                                                                                      -- (terminated)
			csr_readdata      => open,                                                                                     -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                       -- (terminated)
			almost_full_data  => open,                                                                                     -- (terminated)
			almost_empty_data => open,                                                                                     -- (terminated)
			in_empty          => '0',                                                                                      -- (terminated)
			out_empty         => open,                                                                                     -- (terminated)
			in_error          => '0',                                                                                      -- (terminated)
			out_error         => open,                                                                                     -- (terminated)
			in_channel        => '0',                                                                                      -- (terminated)
			out_channel       => open                                                                                      -- (terminated)
		);

	de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 15,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                   --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                            --       clk_reset.reset
			m0_address              => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_src10_ready,                                                                --              cp.ready
			cp_valid                => cmd_xbar_demux_src10_valid,                                                                --                .valid
			cp_data                 => cmd_xbar_demux_src10_data,                                                                 --                .data
			cp_startofpacket        => cmd_xbar_demux_src10_startofpacket,                                                        --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_src10_endofpacket,                                                          --                .endofpacket
			cp_channel              => cmd_xbar_demux_src10_channel,                                                              --                .channel
			rf_sink_ready           => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                      --     (terminated)
			m0_writeresponserequest => open,                                                                                      --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                        --     (terminated)
		);

	de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                   --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			in_data           => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                      -- (terminated)
			csr_read          => '0',                                                                                       -- (terminated)
			csr_write         => '0',                                                                                       -- (terminated)
			csr_readdata      => open,                                                                                      -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                        -- (terminated)
			almost_full_data  => open,                                                                                      -- (terminated)
			almost_empty_data => open,                                                                                      -- (terminated)
			in_empty          => '0',                                                                                       -- (terminated)
			out_empty         => open,                                                                                      -- (terminated)
			in_error          => '0',                                                                                       -- (terminated)
			out_error         => open,                                                                                      -- (terminated)
			in_channel        => '0',                                                                                       -- (terminated)
			out_channel       => open                                                                                       -- (terminated)
		);

	de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 15,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                    --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                             --       clk_reset.reset
			m0_address              => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_src11_ready,                                                                 --              cp.ready
			cp_valid                => cmd_xbar_demux_src11_valid,                                                                 --                .valid
			cp_data                 => cmd_xbar_demux_src11_data,                                                                  --                .data
			cp_startofpacket        => cmd_xbar_demux_src11_startofpacket,                                                         --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_src11_endofpacket,                                                           --                .endofpacket
			cp_channel              => cmd_xbar_demux_src11_channel,                                                               --                .channel
			rf_sink_ready           => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                       --     (terminated)
			m0_writeresponserequest => open,                                                                                       --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                         --     (terminated)
		);

	de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                    --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                             -- clk_reset.reset
			in_data           => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                       -- (terminated)
			csr_read          => '0',                                                                                        -- (terminated)
			csr_write         => '0',                                                                                        -- (terminated)
			csr_readdata      => open,                                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                         -- (terminated)
			almost_full_data  => open,                                                                                       -- (terminated)
			almost_empty_data => open,                                                                                       -- (terminated)
			in_empty          => '0',                                                                                        -- (terminated)
			out_empty         => open,                                                                                       -- (terminated)
			in_error          => '0',                                                                                        -- (terminated)
			out_error         => open,                                                                                       -- (terminated)
			in_channel        => '0',                                                                                        -- (terminated)
			out_channel       => open                                                                                        -- (terminated)
		);

	de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 15,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                   --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                            --       clk_reset.reset
			m0_address              => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_src12_ready,                                                                --              cp.ready
			cp_valid                => cmd_xbar_demux_src12_valid,                                                                --                .valid
			cp_data                 => cmd_xbar_demux_src12_data,                                                                 --                .data
			cp_startofpacket        => cmd_xbar_demux_src12_startofpacket,                                                        --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_src12_endofpacket,                                                          --                .endofpacket
			cp_channel              => cmd_xbar_demux_src12_channel,                                                              --                .channel
			rf_sink_ready           => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                      --     (terminated)
			m0_writeresponserequest => open,                                                                                      --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                        --     (terminated)
		);

	de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2_ht18_lemonde_streit_onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                   --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			in_data           => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                      -- (terminated)
			csr_read          => '0',                                                                                       -- (terminated)
			csr_write         => '0',                                                                                       -- (terminated)
			csr_readdata      => open,                                                                                      -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                        -- (terminated)
			almost_full_data  => open,                                                                                      -- (terminated)
			almost_empty_data => open,                                                                                      -- (terminated)
			in_empty          => '0',                                                                                       -- (terminated)
			out_empty         => open,                                                                                      -- (terminated)
			in_error          => '0',                                                                                       -- (terminated)
			out_error         => open,                                                                                      -- (terminated)
			in_channel        => '0',                                                                                       -- (terminated)
			out_channel       => open                                                                                       -- (terminated)
		);

	sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent : component nios2_ht18_lemonde_streit_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 62,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_ADDR_H                => 42,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 43,
			PKT_TRANS_POSTED          => 44,
			PKT_TRANS_WRITE           => 45,
			PKT_TRANS_READ            => 46,
			PKT_TRANS_LOCK            => 47,
			PKT_SRC_ID_H              => 67,
			PKT_SRC_ID_L              => 64,
			PKT_DEST_ID_H             => 71,
			PKT_DEST_ID_L             => 68,
			PKT_BURSTWRAP_H           => 54,
			PKT_BURSTWRAP_L           => 52,
			PKT_BYTE_CNT_H            => 51,
			PKT_BYTE_CNT_L            => 49,
			PKT_PROTECTION_H          => 75,
			PKT_PROTECTION_L          => 73,
			PKT_RESPONSE_STATUS_H     => 81,
			PKT_RESPONSE_STATUS_L     => 80,
			PKT_BURST_SIZE_H          => 57,
			PKT_BURST_SIZE_L          => 55,
			ST_CHANNEL_W              => 15,
			ST_DATA_W                 => 82,
			AVS_BURSTCOUNT_W          => 2,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                     --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                              --       clk_reset.reset
			m0_address              => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_source0_ready,                                                                 --              cp.ready
			cp_valid                => burst_adapter_source0_valid,                                                                 --                .valid
			cp_data                 => burst_adapter_source0_data,                                                                  --                .data
			cp_startofpacket        => burst_adapter_source0_startofpacket,                                                         --                .startofpacket
			cp_endofpacket          => burst_adapter_source0_endofpacket,                                                           --                .endofpacket
			cp_channel              => burst_adapter_source0_channel,                                                               --                .channel
			rf_sink_ready           => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                          --     (terminated)
		);

	sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2_ht18_lemonde_streit_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 83,
			FIFO_DEPTH          => 3,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                     --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                              -- clk_reset.reset
			in_data           => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                        -- (terminated)
			csr_read          => '0',                                                                                         -- (terminated)
			csr_write         => '0',                                                                                         -- (terminated)
			csr_readdata      => open,                                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                          -- (terminated)
			almost_full_data  => open,                                                                                        -- (terminated)
			almost_empty_data => open,                                                                                        -- (terminated)
			in_empty          => '0',                                                                                         -- (terminated)
			out_empty         => open,                                                                                        -- (terminated)
			in_error          => '0',                                                                                         -- (terminated)
			out_error         => open,                                                                                        -- (terminated)
			in_channel        => '0',                                                                                         -- (terminated)
			out_channel       => open                                                                                         -- (terminated)
		);

	sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2_ht18_lemonde_streit_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 18,
			FIFO_DEPTH          => 3,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                               --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			in_data           => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                                  -- (terminated)
			csr_read          => '0',                                                                                   -- (terminated)
			csr_write         => '0',                                                                                   -- (terminated)
			csr_readdata      => open,                                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                    -- (terminated)
			almost_full_data  => open,                                                                                  -- (terminated)
			almost_empty_data => open,                                                                                  -- (terminated)
			in_startofpacket  => '0',                                                                                   -- (terminated)
			in_endofpacket    => '0',                                                                                   -- (terminated)
			out_startofpacket => open,                                                                                  -- (terminated)
			out_endofpacket   => open,                                                                                  -- (terminated)
			in_empty          => '0',                                                                                   -- (terminated)
			out_empty         => open,                                                                                  -- (terminated)
			in_error          => '0',                                                                                   -- (terminated)
			out_error         => open,                                                                                  -- (terminated)
			in_channel        => '0',                                                                                   -- (terminated)
			out_channel       => open                                                                                   -- (terminated)
		);

	sdram_s1_translator_avalon_universal_slave_0_agent : component nios2_ht18_lemonde_streit_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 62,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_ADDR_H                => 42,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 43,
			PKT_TRANS_POSTED          => 44,
			PKT_TRANS_WRITE           => 45,
			PKT_TRANS_READ            => 46,
			PKT_TRANS_LOCK            => 47,
			PKT_SRC_ID_H              => 67,
			PKT_SRC_ID_L              => 64,
			PKT_DEST_ID_H             => 71,
			PKT_DEST_ID_L             => 68,
			PKT_BURSTWRAP_H           => 54,
			PKT_BURSTWRAP_L           => 52,
			PKT_BYTE_CNT_H            => 51,
			PKT_BYTE_CNT_L            => 49,
			PKT_PROTECTION_H          => 75,
			PKT_PROTECTION_L          => 73,
			PKT_RESPONSE_STATUS_H     => 81,
			PKT_RESPONSE_STATUS_L     => 80,
			PKT_BURST_SIZE_H          => 57,
			PKT_BURST_SIZE_L          => 55,
			ST_CHANNEL_W              => 15,
			ST_DATA_W                 => 82,
			AVS_BURSTCOUNT_W          => 2,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                       --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                --       clk_reset.reset
			m0_address              => sdram_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sdram_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sdram_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sdram_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_001_source0_ready,                                               --              cp.ready
			cp_valid                => burst_adapter_001_source0_valid,                                               --                .valid
			cp_data                 => burst_adapter_001_source0_data,                                                --                .data
			cp_startofpacket        => burst_adapter_001_source0_startofpacket,                                       --                .startofpacket
			cp_endofpacket          => burst_adapter_001_source0_endofpacket,                                         --                .endofpacket
			cp_channel              => burst_adapter_001_source0_channel,                                             --                .channel
			rf_sink_ready           => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                          --     (terminated)
			m0_writeresponserequest => open,                                                                          --     (terminated)
			m0_writeresponsevalid   => '0'                                                                            --     (terminated)
		);

	sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2_ht18_lemonde_streit_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 83,
			FIFO_DEPTH          => 8,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                       --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                -- clk_reset.reset
			in_data           => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                          -- (terminated)
			csr_read          => '0',                                                                           -- (terminated)
			csr_write         => '0',                                                                           -- (terminated)
			csr_readdata      => open,                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                            -- (terminated)
			almost_full_data  => open,                                                                          -- (terminated)
			almost_empty_data => open,                                                                          -- (terminated)
			in_empty          => '0',                                                                           -- (terminated)
			out_empty         => open,                                                                          -- (terminated)
			in_error          => '0',                                                                           -- (terminated)
			out_error         => open,                                                                          -- (terminated)
			in_channel        => '0',                                                                           -- (terminated)
			out_channel       => open                                                                           -- (terminated)
		);

	sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2_ht18_lemonde_streit_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 18,
			FIFO_DEPTH          => 8,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 3,
			USE_MEMORY_BLOCKS   => 1,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                 --       clk.clk
			reset             => rst_controller_reset_out_reset,                                          -- clk_reset.reset
			in_data           => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                    -- (terminated)
			csr_read          => '0',                                                                     -- (terminated)
			csr_write         => '0',                                                                     -- (terminated)
			csr_readdata      => open,                                                                    -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                      -- (terminated)
			almost_full_data  => open,                                                                    -- (terminated)
			almost_empty_data => open,                                                                    -- (terminated)
			in_startofpacket  => '0',                                                                     -- (terminated)
			in_endofpacket    => '0',                                                                     -- (terminated)
			out_startofpacket => open,                                                                    -- (terminated)
			out_endofpacket   => open,                                                                    -- (terminated)
			in_empty          => '0',                                                                     -- (terminated)
			out_empty         => open,                                                                    -- (terminated)
			in_error          => '0',                                                                     -- (terminated)
			out_error         => open,                                                                    -- (terminated)
			in_channel        => '0',                                                                     -- (terminated)
			out_channel       => open                                                                     -- (terminated)
		);

	addr_router : component nios2_ht18_lemonde_streit_addr_router
		port map (
			sink_ready         => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_ht18_lemonde_streit_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                                           --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                                    -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                                             --       src.ready
			src_valid          => addr_router_src_valid,                                                                             --          .valid
			src_data           => addr_router_src_data,                                                                              --          .data
			src_channel        => addr_router_src_channel,                                                                           --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                                     --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                                        --          .endofpacket
		);

	addr_router_001 : component nios2_ht18_lemonde_streit_addr_router_001
		port map (
			sink_ready         => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_ht18_lemonde_streit_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                                           -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                                                --       src.ready
			src_valid          => addr_router_001_src_valid,                                                                                --          .valid
			src_data           => addr_router_001_src_data,                                                                                 --          .data
			src_channel        => addr_router_001_src_channel,                                                                              --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                                                        --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                                                           --          .endofpacket
		);

	id_router : component nios2_ht18_lemonde_streit_id_router
		port map (
			sink_ready         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                         --       src.ready
			src_valid          => id_router_src_valid,                                                         --          .valid
			src_data           => id_router_src_data,                                                          --          .data
			src_channel        => id_router_src_channel,                                                       --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                 --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                    --          .endofpacket
		);

	id_router_001 : component nios2_ht18_lemonde_streit_id_router_001
		port map (
			sink_ready         => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => ht18_lemonde_streit_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                                      --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                           -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                                                      --       src.ready
			src_valid          => id_router_001_src_valid,                                                                      --          .valid
			src_data           => id_router_001_src_data,                                                                       --          .data
			src_channel        => id_router_001_src_channel,                                                                    --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                                              --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                                                 --          .endofpacket
		);

	id_router_002 : component nios2_ht18_lemonde_streit_id_router_001
		port map (
			sink_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                           -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                                                  --       src.ready
			src_valid          => id_router_002_src_valid,                                                                  --          .valid
			src_data           => id_router_002_src_data,                                                                   --          .data
			src_channel        => id_router_002_src_channel,                                                                --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                                          --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                                             --          .endofpacket
		);

	id_router_003 : component nios2_ht18_lemonde_streit_id_router
		port map (
			sink_ready         => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_ht18_lemonde_streit_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                                                --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                                         -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                                                                --       src.ready
			src_valid          => id_router_003_src_valid,                                                                                --          .valid
			src_data           => id_router_003_src_data,                                                                                 --          .data
			src_channel        => id_router_003_src_channel,                                                                              --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                                                        --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                                                           --          .endofpacket
		);

	id_router_004 : component nios2_ht18_lemonde_streit_id_router_001
		port map (
			sink_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                               --       src.ready
			src_valid          => id_router_004_src_valid,                                               --          .valid
			src_data           => id_router_004_src_data,                                                --          .data
			src_channel        => id_router_004_src_channel,                                             --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                          --          .endofpacket
		);

	id_router_005 : component nios2_ht18_lemonde_streit_id_router_001
		port map (
			sink_ready         => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                               --       src.ready
			src_valid          => id_router_005_src_valid,                                               --          .valid
			src_data           => id_router_005_src_data,                                                --          .data
			src_channel        => id_router_005_src_channel,                                             --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                          --          .endofpacket
		);

	id_router_006 : component nios2_ht18_lemonde_streit_id_router_001
		port map (
			sink_ready         => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => p_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                                            --       src.ready
			src_valid          => id_router_006_src_valid,                                                            --          .valid
			src_data           => id_router_006_src_data,                                                             --          .data
			src_channel        => id_router_006_src_channel,                                                          --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                                    --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                                       --          .endofpacket
		);

	id_router_007 : component nios2_ht18_lemonde_streit_id_router_001
		port map (
			sink_ready         => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => de2_pio_toggles18_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                         --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			src_ready          => id_router_007_src_ready,                                                         --       src.ready
			src_valid          => id_router_007_src_valid,                                                         --          .valid
			src_data           => id_router_007_src_data,                                                          --          .data
			src_channel        => id_router_007_src_channel,                                                       --          .channel
			src_startofpacket  => id_router_007_src_startofpacket,                                                 --          .startofpacket
			src_endofpacket    => id_router_007_src_endofpacket                                                    --          .endofpacket
		);

	id_router_008 : component nios2_ht18_lemonde_streit_id_router_001
		port map (
			sink_ready         => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => de2_pio_keys4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => id_router_008_src_ready,                                                     --       src.ready
			src_valid          => id_router_008_src_valid,                                                     --          .valid
			src_data           => id_router_008_src_data,                                                      --          .data
			src_channel        => id_router_008_src_channel,                                                   --          .channel
			src_startofpacket  => id_router_008_src_startofpacket,                                             --          .startofpacket
			src_endofpacket    => id_router_008_src_endofpacket                                                --          .endofpacket
		);

	id_router_009 : component nios2_ht18_lemonde_streit_id_router_001
		port map (
			sink_ready         => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => de2_pio_redled18_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                        --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                 -- clk_reset.reset
			src_ready          => id_router_009_src_ready,                                                        --       src.ready
			src_valid          => id_router_009_src_valid,                                                        --          .valid
			src_data           => id_router_009_src_data,                                                         --          .data
			src_channel        => id_router_009_src_channel,                                                      --          .channel
			src_startofpacket  => id_router_009_src_startofpacket,                                                --          .startofpacket
			src_endofpacket    => id_router_009_src_endofpacket                                                   --          .endofpacket
		);

	id_router_010 : component nios2_ht18_lemonde_streit_id_router_001
		port map (
			sink_ready         => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => de2_pio_greenled9_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                         --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			src_ready          => id_router_010_src_ready,                                                         --       src.ready
			src_valid          => id_router_010_src_valid,                                                         --          .valid
			src_data           => id_router_010_src_data,                                                          --          .data
			src_channel        => id_router_010_src_channel,                                                       --          .channel
			src_startofpacket  => id_router_010_src_startofpacket,                                                 --          .startofpacket
			src_endofpacket    => id_router_010_src_endofpacket                                                    --          .endofpacket
		);

	id_router_011 : component nios2_ht18_lemonde_streit_id_router_001
		port map (
			sink_ready         => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => de2_pio_hex_high28_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                          --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			src_ready          => id_router_011_src_ready,                                                          --       src.ready
			src_valid          => id_router_011_src_valid,                                                          --          .valid
			src_data           => id_router_011_src_data,                                                           --          .data
			src_channel        => id_router_011_src_channel,                                                        --          .channel
			src_startofpacket  => id_router_011_src_startofpacket,                                                  --          .startofpacket
			src_endofpacket    => id_router_011_src_endofpacket                                                     --          .endofpacket
		);

	id_router_012 : component nios2_ht18_lemonde_streit_id_router_001
		port map (
			sink_ready         => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => de2_pio_hex_low28_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                         --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			src_ready          => id_router_012_src_ready,                                                         --       src.ready
			src_valid          => id_router_012_src_valid,                                                         --          .valid
			src_data           => id_router_012_src_data,                                                          --          .data
			src_channel        => id_router_012_src_channel,                                                       --          .channel
			src_startofpacket  => id_router_012_src_startofpacket,                                                 --          .startofpacket
			src_endofpacket    => id_router_012_src_endofpacket                                                    --          .endofpacket
		);

	id_router_013 : component nios2_ht18_lemonde_streit_id_router_013
		port map (
			sink_ready         => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                           --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                    -- clk_reset.reset
			src_ready          => id_router_013_src_ready,                                                           --       src.ready
			src_valid          => id_router_013_src_valid,                                                           --          .valid
			src_data           => id_router_013_src_data,                                                            --          .data
			src_channel        => id_router_013_src_channel,                                                         --          .channel
			src_startofpacket  => id_router_013_src_startofpacket,                                                   --          .startofpacket
			src_endofpacket    => id_router_013_src_endofpacket                                                      --          .endofpacket
		);

	id_router_014 : component nios2_ht18_lemonde_streit_id_router_013
		port map (
			sink_ready         => sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sdram_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                             --       clk.clk
			reset              => rst_controller_reset_out_reset,                                      -- clk_reset.reset
			src_ready          => id_router_014_src_ready,                                             --       src.ready
			src_valid          => id_router_014_src_valid,                                             --          .valid
			src_data           => id_router_014_src_data,                                              --          .data
			src_channel        => id_router_014_src_channel,                                           --          .channel
			src_startofpacket  => id_router_014_src_startofpacket,                                     --          .startofpacket
			src_endofpacket    => id_router_014_src_endofpacket                                        --          .endofpacket
		);

	burst_adapter : component altera_merlin_burst_adapter
		generic map (
			PKT_ADDR_H                => 42,
			PKT_ADDR_L                => 18,
			PKT_BEGIN_BURST           => 62,
			PKT_BYTE_CNT_H            => 51,
			PKT_BYTE_CNT_L            => 49,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_BURST_SIZE_H          => 57,
			PKT_BURST_SIZE_L          => 55,
			PKT_BURST_TYPE_H          => 59,
			PKT_BURST_TYPE_L          => 58,
			PKT_BURSTWRAP_H           => 54,
			PKT_BURSTWRAP_L           => 52,
			PKT_TRANS_COMPRESSED_READ => 43,
			PKT_TRANS_WRITE           => 45,
			PKT_TRANS_READ            => 46,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 82,
			ST_CHANNEL_W              => 15,
			OUT_BYTE_CNT_H            => 50,
			OUT_BURSTWRAP_H           => 54,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 3,
			BURSTWRAP_CONST_VALUE     => 3
		)
		port map (
			clk                   => up_clocks_0_sys_clk_clk,             --       cr0.clk
			reset                 => rst_controller_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => width_adapter_src_valid,             --     sink0.valid
			sink0_data            => width_adapter_src_data,              --          .data
			sink0_channel         => width_adapter_src_channel,           --          .channel
			sink0_startofpacket   => width_adapter_src_startofpacket,     --          .startofpacket
			sink0_endofpacket     => width_adapter_src_endofpacket,       --          .endofpacket
			sink0_ready           => width_adapter_src_ready,             --          .ready
			source0_valid         => burst_adapter_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_source0_data,          --          .data
			source0_channel       => burst_adapter_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_source0_ready          --          .ready
		);

	burst_adapter_001 : component altera_merlin_burst_adapter
		generic map (
			PKT_ADDR_H                => 42,
			PKT_ADDR_L                => 18,
			PKT_BEGIN_BURST           => 62,
			PKT_BYTE_CNT_H            => 51,
			PKT_BYTE_CNT_L            => 49,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_BURST_SIZE_H          => 57,
			PKT_BURST_SIZE_L          => 55,
			PKT_BURST_TYPE_H          => 59,
			PKT_BURST_TYPE_L          => 58,
			PKT_BURSTWRAP_H           => 54,
			PKT_BURSTWRAP_L           => 52,
			PKT_TRANS_COMPRESSED_READ => 43,
			PKT_TRANS_WRITE           => 45,
			PKT_TRANS_READ            => 46,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 82,
			ST_CHANNEL_W              => 15,
			OUT_BYTE_CNT_H            => 50,
			OUT_BURSTWRAP_H           => 54,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 3,
			BURSTWRAP_CONST_VALUE     => 3
		)
		port map (
			clk                   => up_clocks_0_sys_clk_clk,                 --       cr0.clk
			reset                 => rst_controller_reset_out_reset,          -- cr0_reset.reset
			sink0_valid           => width_adapter_002_src_valid,             --     sink0.valid
			sink0_data            => width_adapter_002_src_data,              --          .data
			sink0_channel         => width_adapter_002_src_channel,           --          .channel
			sink0_startofpacket   => width_adapter_002_src_startofpacket,     --          .startofpacket
			sink0_endofpacket     => width_adapter_002_src_endofpacket,       --          .endofpacket
			sink0_ready           => width_adapter_002_src_ready,             --          .ready
			source0_valid         => burst_adapter_001_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_001_source0_data,          --          .data
			source0_channel       => burst_adapter_001_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_001_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_001_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_001_source0_ready          --          .ready
		);

	rst_controller : component nios2_ht18_lemonde_streit_rst_controller
		generic map (
			NUM_RESET_INPUTS        => 2,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 1
		)
		port map (
			reset_in0  => nios2_ht18_lemonde_streit_jtag_debug_module_reset_reset, -- reset_in0.reset
			reset_in1  => reset_reset_n_ports_inv,                                 -- reset_in1.reset
			clk        => up_clocks_0_sys_clk_clk,                                 --       clk.clk
			reset_out  => rst_controller_reset_out_reset,                          -- reset_out.reset
			reset_req  => rst_controller_reset_out_reset_req,                      --          .reset_req
			reset_in2  => '0',                                                     -- (terminated)
			reset_in3  => '0',                                                     -- (terminated)
			reset_in4  => '0',                                                     -- (terminated)
			reset_in5  => '0',                                                     -- (terminated)
			reset_in6  => '0',                                                     -- (terminated)
			reset_in7  => '0',                                                     -- (terminated)
			reset_in8  => '0',                                                     -- (terminated)
			reset_in9  => '0',                                                     -- (terminated)
			reset_in10 => '0',                                                     -- (terminated)
			reset_in11 => '0',                                                     -- (terminated)
			reset_in12 => '0',                                                     -- (terminated)
			reset_in13 => '0',                                                     -- (terminated)
			reset_in14 => '0',                                                     -- (terminated)
			reset_in15 => '0'                                                      -- (terminated)
		);

	rst_controller_001 : component nios2_ht18_lemonde_streit_rst_controller_001
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk        => up_clocks_0_sys_clk_clk,            --       clk.clk
			reset_out  => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req  => open,                               -- (terminated)
			reset_in1  => '0',                                -- (terminated)
			reset_in2  => '0',                                -- (terminated)
			reset_in3  => '0',                                -- (terminated)
			reset_in4  => '0',                                -- (terminated)
			reset_in5  => '0',                                -- (terminated)
			reset_in6  => '0',                                -- (terminated)
			reset_in7  => '0',                                -- (terminated)
			reset_in8  => '0',                                -- (terminated)
			reset_in9  => '0',                                -- (terminated)
			reset_in10 => '0',                                -- (terminated)
			reset_in11 => '0',                                -- (terminated)
			reset_in12 => '0',                                -- (terminated)
			reset_in13 => '0',                                -- (terminated)
			reset_in14 => '0',                                -- (terminated)
			reset_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component nios2_ht18_lemonde_streit_rst_controller_002
		generic map (
			NUM_RESET_INPUTS        => 2,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,                                 -- reset_in0.reset
			reset_in1  => nios2_ht18_lemonde_streit_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk        => clk_clk,                                                 --       clk.clk
			reset_out  => rst_controller_002_reset_out_reset,                      -- reset_out.reset
			reset_req  => open,                                                    -- (terminated)
			reset_in2  => '0',                                                     -- (terminated)
			reset_in3  => '0',                                                     -- (terminated)
			reset_in4  => '0',                                                     -- (terminated)
			reset_in5  => '0',                                                     -- (terminated)
			reset_in6  => '0',                                                     -- (terminated)
			reset_in7  => '0',                                                     -- (terminated)
			reset_in8  => '0',                                                     -- (terminated)
			reset_in9  => '0',                                                     -- (terminated)
			reset_in10 => '0',                                                     -- (terminated)
			reset_in11 => '0',                                                     -- (terminated)
			reset_in12 => '0',                                                     -- (terminated)
			reset_in13 => '0',                                                     -- (terminated)
			reset_in14 => '0',                                                     -- (terminated)
			reset_in15 => '0'                                                      -- (terminated)
		);

	cmd_xbar_demux : component nios2_ht18_lemonde_streit_cmd_xbar_demux
		port map (
			clk                 => up_clocks_0_sys_clk_clk,            --       clk.clk
			reset               => rst_controller_reset_out_reset,     -- clk_reset.reset
			sink_ready          => addr_router_src_ready,              --      sink.ready
			sink_channel        => addr_router_src_channel,            --          .channel
			sink_data           => addr_router_src_data,               --          .data
			sink_startofpacket  => addr_router_src_startofpacket,      --          .startofpacket
			sink_endofpacket    => addr_router_src_endofpacket,        --          .endofpacket
			sink_valid(0)       => addr_router_src_valid,              --          .valid
			src0_ready          => cmd_xbar_demux_src0_ready,          --      src0.ready
			src0_valid          => cmd_xbar_demux_src0_valid,          --          .valid
			src0_data           => cmd_xbar_demux_src0_data,           --          .data
			src0_channel        => cmd_xbar_demux_src0_channel,        --          .channel
			src0_startofpacket  => cmd_xbar_demux_src0_startofpacket,  --          .startofpacket
			src0_endofpacket    => cmd_xbar_demux_src0_endofpacket,    --          .endofpacket
			src1_ready          => cmd_xbar_demux_src1_ready,          --      src1.ready
			src1_valid          => cmd_xbar_demux_src1_valid,          --          .valid
			src1_data           => cmd_xbar_demux_src1_data,           --          .data
			src1_channel        => cmd_xbar_demux_src1_channel,        --          .channel
			src1_startofpacket  => cmd_xbar_demux_src1_startofpacket,  --          .startofpacket
			src1_endofpacket    => cmd_xbar_demux_src1_endofpacket,    --          .endofpacket
			src2_ready          => cmd_xbar_demux_src2_ready,          --      src2.ready
			src2_valid          => cmd_xbar_demux_src2_valid,          --          .valid
			src2_data           => cmd_xbar_demux_src2_data,           --          .data
			src2_channel        => cmd_xbar_demux_src2_channel,        --          .channel
			src2_startofpacket  => cmd_xbar_demux_src2_startofpacket,  --          .startofpacket
			src2_endofpacket    => cmd_xbar_demux_src2_endofpacket,    --          .endofpacket
			src3_ready          => cmd_xbar_demux_src3_ready,          --      src3.ready
			src3_valid          => cmd_xbar_demux_src3_valid,          --          .valid
			src3_data           => cmd_xbar_demux_src3_data,           --          .data
			src3_channel        => cmd_xbar_demux_src3_channel,        --          .channel
			src3_startofpacket  => cmd_xbar_demux_src3_startofpacket,  --          .startofpacket
			src3_endofpacket    => cmd_xbar_demux_src3_endofpacket,    --          .endofpacket
			src4_ready          => cmd_xbar_demux_src4_ready,          --      src4.ready
			src4_valid          => cmd_xbar_demux_src4_valid,          --          .valid
			src4_data           => cmd_xbar_demux_src4_data,           --          .data
			src4_channel        => cmd_xbar_demux_src4_channel,        --          .channel
			src4_startofpacket  => cmd_xbar_demux_src4_startofpacket,  --          .startofpacket
			src4_endofpacket    => cmd_xbar_demux_src4_endofpacket,    --          .endofpacket
			src5_ready          => cmd_xbar_demux_src5_ready,          --      src5.ready
			src5_valid          => cmd_xbar_demux_src5_valid,          --          .valid
			src5_data           => cmd_xbar_demux_src5_data,           --          .data
			src5_channel        => cmd_xbar_demux_src5_channel,        --          .channel
			src5_startofpacket  => cmd_xbar_demux_src5_startofpacket,  --          .startofpacket
			src5_endofpacket    => cmd_xbar_demux_src5_endofpacket,    --          .endofpacket
			src6_ready          => cmd_xbar_demux_src6_ready,          --      src6.ready
			src6_valid          => cmd_xbar_demux_src6_valid,          --          .valid
			src6_data           => cmd_xbar_demux_src6_data,           --          .data
			src6_channel        => cmd_xbar_demux_src6_channel,        --          .channel
			src6_startofpacket  => cmd_xbar_demux_src6_startofpacket,  --          .startofpacket
			src6_endofpacket    => cmd_xbar_demux_src6_endofpacket,    --          .endofpacket
			src7_ready          => cmd_xbar_demux_src7_ready,          --      src7.ready
			src7_valid          => cmd_xbar_demux_src7_valid,          --          .valid
			src7_data           => cmd_xbar_demux_src7_data,           --          .data
			src7_channel        => cmd_xbar_demux_src7_channel,        --          .channel
			src7_startofpacket  => cmd_xbar_demux_src7_startofpacket,  --          .startofpacket
			src7_endofpacket    => cmd_xbar_demux_src7_endofpacket,    --          .endofpacket
			src8_ready          => cmd_xbar_demux_src8_ready,          --      src8.ready
			src8_valid          => cmd_xbar_demux_src8_valid,          --          .valid
			src8_data           => cmd_xbar_demux_src8_data,           --          .data
			src8_channel        => cmd_xbar_demux_src8_channel,        --          .channel
			src8_startofpacket  => cmd_xbar_demux_src8_startofpacket,  --          .startofpacket
			src8_endofpacket    => cmd_xbar_demux_src8_endofpacket,    --          .endofpacket
			src9_ready          => cmd_xbar_demux_src9_ready,          --      src9.ready
			src9_valid          => cmd_xbar_demux_src9_valid,          --          .valid
			src9_data           => cmd_xbar_demux_src9_data,           --          .data
			src9_channel        => cmd_xbar_demux_src9_channel,        --          .channel
			src9_startofpacket  => cmd_xbar_demux_src9_startofpacket,  --          .startofpacket
			src9_endofpacket    => cmd_xbar_demux_src9_endofpacket,    --          .endofpacket
			src10_ready         => cmd_xbar_demux_src10_ready,         --     src10.ready
			src10_valid         => cmd_xbar_demux_src10_valid,         --          .valid
			src10_data          => cmd_xbar_demux_src10_data,          --          .data
			src10_channel       => cmd_xbar_demux_src10_channel,       --          .channel
			src10_startofpacket => cmd_xbar_demux_src10_startofpacket, --          .startofpacket
			src10_endofpacket   => cmd_xbar_demux_src10_endofpacket,   --          .endofpacket
			src11_ready         => cmd_xbar_demux_src11_ready,         --     src11.ready
			src11_valid         => cmd_xbar_demux_src11_valid,         --          .valid
			src11_data          => cmd_xbar_demux_src11_data,          --          .data
			src11_channel       => cmd_xbar_demux_src11_channel,       --          .channel
			src11_startofpacket => cmd_xbar_demux_src11_startofpacket, --          .startofpacket
			src11_endofpacket   => cmd_xbar_demux_src11_endofpacket,   --          .endofpacket
			src12_ready         => cmd_xbar_demux_src12_ready,         --     src12.ready
			src12_valid         => cmd_xbar_demux_src12_valid,         --          .valid
			src12_data          => cmd_xbar_demux_src12_data,          --          .data
			src12_channel       => cmd_xbar_demux_src12_channel,       --          .channel
			src12_startofpacket => cmd_xbar_demux_src12_startofpacket, --          .startofpacket
			src12_endofpacket   => cmd_xbar_demux_src12_endofpacket,   --          .endofpacket
			src13_ready         => cmd_xbar_demux_src13_ready,         --     src13.ready
			src13_valid         => cmd_xbar_demux_src13_valid,         --          .valid
			src13_data          => cmd_xbar_demux_src13_data,          --          .data
			src13_channel       => cmd_xbar_demux_src13_channel,       --          .channel
			src13_startofpacket => cmd_xbar_demux_src13_startofpacket, --          .startofpacket
			src13_endofpacket   => cmd_xbar_demux_src13_endofpacket,   --          .endofpacket
			src14_ready         => cmd_xbar_demux_src14_ready,         --     src14.ready
			src14_valid         => cmd_xbar_demux_src14_valid,         --          .valid
			src14_data          => cmd_xbar_demux_src14_data,          --          .data
			src14_channel       => cmd_xbar_demux_src14_channel,       --          .channel
			src14_startofpacket => cmd_xbar_demux_src14_startofpacket, --          .startofpacket
			src14_endofpacket   => cmd_xbar_demux_src14_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_001 : component nios2_ht18_lemonde_streit_cmd_xbar_demux_001
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_001_src_ready,             --      sink.ready
			sink_channel       => addr_router_001_src_channel,           --          .channel
			sink_data          => addr_router_001_src_data,              --          .data
			sink_startofpacket => addr_router_001_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_001_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_001_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_001_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => cmd_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			src1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			src2_ready         => cmd_xbar_demux_001_src2_ready,         --      src2.ready
			src2_valid         => cmd_xbar_demux_001_src2_valid,         --          .valid
			src2_data          => cmd_xbar_demux_001_src2_data,          --          .data
			src2_channel       => cmd_xbar_demux_001_src2_channel,       --          .channel
			src2_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --          .startofpacket
			src2_endofpacket   => cmd_xbar_demux_001_src2_endofpacket,   --          .endofpacket
			src3_ready         => cmd_xbar_demux_001_src3_ready,         --      src3.ready
			src3_valid         => cmd_xbar_demux_001_src3_valid,         --          .valid
			src3_data          => cmd_xbar_demux_001_src3_data,          --          .data
			src3_channel       => cmd_xbar_demux_001_src3_channel,       --          .channel
			src3_startofpacket => cmd_xbar_demux_001_src3_startofpacket, --          .startofpacket
			src3_endofpacket   => cmd_xbar_demux_001_src3_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux : component nios2_ht18_lemonde_streit_cmd_xbar_mux
		port map (
			clk                 => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_003 : component nios2_ht18_lemonde_streit_cmd_xbar_mux
		port map (
			clk                 => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_003_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_003_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_003_src_data,             --          .data
			src_channel         => cmd_xbar_mux_003_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_003_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_003_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src3_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src3_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src3_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src3_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src3_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src3_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_013 : component nios2_ht18_lemonde_streit_cmd_xbar_mux
		port map (
			clk                 => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_013_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_013_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_013_src_data,             --          .data
			src_channel         => cmd_xbar_mux_013_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_013_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_013_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src13_ready,            --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src13_valid,            --          .valid
			sink0_channel       => cmd_xbar_demux_src13_channel,          --          .channel
			sink0_data          => cmd_xbar_demux_src13_data,             --          .data
			sink0_startofpacket => cmd_xbar_demux_src13_startofpacket,    --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src13_endofpacket,      --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src2_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src2_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src2_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src2_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src2_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_014 : component nios2_ht18_lemonde_streit_cmd_xbar_mux
		port map (
			clk                 => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_014_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_014_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_014_src_data,             --          .data
			src_channel         => cmd_xbar_mux_014_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_014_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_014_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src14_ready,            --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src14_valid,            --          .valid
			sink0_channel       => cmd_xbar_demux_src14_channel,          --          .channel
			sink0_data          => cmd_xbar_demux_src14_data,             --          .data
			sink0_startofpacket => cmd_xbar_demux_src14_startofpacket,    --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src14_endofpacket,      --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src3_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src3_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src3_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src3_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src3_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src3_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux : component nios2_ht18_lemonde_streit_rsp_xbar_demux
		port map (
			clk                => up_clocks_0_sys_clk_clk,           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_src_ready,               --      sink.ready
			sink_channel       => id_router_src_channel,             --          .channel
			sink_data          => id_router_src_data,                --          .data
			sink_startofpacket => id_router_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_001 : component nios2_ht18_lemonde_streit_rsp_xbar_demux_001
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_001_src_ready,               --      sink.ready
			sink_channel       => id_router_001_src_channel,             --          .channel
			sink_data          => id_router_001_src_data,                --          .data
			sink_startofpacket => id_router_001_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_001_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_001_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component nios2_ht18_lemonde_streit_rsp_xbar_demux_001
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_002_src_ready,               --      sink.ready
			sink_channel       => id_router_002_src_channel,             --          .channel
			sink_data          => id_router_002_src_data,                --          .data
			sink_startofpacket => id_router_002_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_002_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_002_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component nios2_ht18_lemonde_streit_rsp_xbar_demux
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_003_src_ready,               --      sink.ready
			sink_channel       => id_router_003_src_channel,             --          .channel
			sink_data          => id_router_003_src_data,                --          .data
			sink_startofpacket => id_router_003_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_003_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_003_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_003_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_003_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_003_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_003_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_003_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_004 : component nios2_ht18_lemonde_streit_rsp_xbar_demux_001
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_004_src_ready,               --      sink.ready
			sink_channel       => id_router_004_src_channel,             --          .channel
			sink_data          => id_router_004_src_data,                --          .data
			sink_startofpacket => id_router_004_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_004_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_004_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_005 : component nios2_ht18_lemonde_streit_rsp_xbar_demux_001
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_005_src_ready,               --      sink.ready
			sink_channel       => id_router_005_src_channel,             --          .channel
			sink_data          => id_router_005_src_data,                --          .data
			sink_startofpacket => id_router_005_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_005_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_005_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_006 : component nios2_ht18_lemonde_streit_rsp_xbar_demux_001
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_006_src_ready,               --      sink.ready
			sink_channel       => id_router_006_src_channel,             --          .channel
			sink_data          => id_router_006_src_data,                --          .data
			sink_startofpacket => id_router_006_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_006_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_006_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_007 : component nios2_ht18_lemonde_streit_rsp_xbar_demux_001
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_007_src_ready,               --      sink.ready
			sink_channel       => id_router_007_src_channel,             --          .channel
			sink_data          => id_router_007_src_data,                --          .data
			sink_startofpacket => id_router_007_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_007_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_007_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_007_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_007_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_007_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_008 : component nios2_ht18_lemonde_streit_rsp_xbar_demux_001
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_008_src_ready,               --      sink.ready
			sink_channel       => id_router_008_src_channel,             --          .channel
			sink_data          => id_router_008_src_data,                --          .data
			sink_startofpacket => id_router_008_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_008_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_008_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_008_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_008_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_008_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_009 : component nios2_ht18_lemonde_streit_rsp_xbar_demux_001
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_009_src_ready,               --      sink.ready
			sink_channel       => id_router_009_src_channel,             --          .channel
			sink_data          => id_router_009_src_data,                --          .data
			sink_startofpacket => id_router_009_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_009_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_009_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_009_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_009_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_009_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_010 : component nios2_ht18_lemonde_streit_rsp_xbar_demux_001
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_010_src_ready,               --      sink.ready
			sink_channel       => id_router_010_src_channel,             --          .channel
			sink_data          => id_router_010_src_data,                --          .data
			sink_startofpacket => id_router_010_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_010_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_010_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_010_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_010_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_010_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_011 : component nios2_ht18_lemonde_streit_rsp_xbar_demux_001
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_011_src_ready,               --      sink.ready
			sink_channel       => id_router_011_src_channel,             --          .channel
			sink_data          => id_router_011_src_data,                --          .data
			sink_startofpacket => id_router_011_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_011_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_011_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_011_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_011_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_011_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_012 : component nios2_ht18_lemonde_streit_rsp_xbar_demux_001
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_012_src_ready,               --      sink.ready
			sink_channel       => id_router_012_src_channel,             --          .channel
			sink_data          => id_router_012_src_data,                --          .data
			sink_startofpacket => id_router_012_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_012_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_012_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_012_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_012_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_012_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_013 : component nios2_ht18_lemonde_streit_rsp_xbar_demux
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => width_adapter_001_src_ready,           --      sink.ready
			sink_channel       => width_adapter_001_src_channel,         --          .channel
			sink_data          => width_adapter_001_src_data,            --          .data
			sink_startofpacket => width_adapter_001_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_001_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_001_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_013_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_013_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_013_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_013_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_013_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_013_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_013_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_013_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_013_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_014 : component nios2_ht18_lemonde_streit_rsp_xbar_demux
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => width_adapter_003_src_ready,           --      sink.ready
			sink_channel       => width_adapter_003_src_channel,         --          .channel
			sink_data          => width_adapter_003_src_data,            --          .data
			sink_startofpacket => width_adapter_003_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_003_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_003_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_014_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_014_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_014_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_014_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_014_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_014_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_014_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_014_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_014_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_014_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_014_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_014_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component nios2_ht18_lemonde_streit_rsp_xbar_mux
		port map (
			clk                  => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready            => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid            => rsp_xbar_mux_src_valid,                --          .valid
			src_data             => rsp_xbar_mux_src_data,                 --          .data
			src_channel          => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket    => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket      => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready          => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid          => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel        => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data           => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket  => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket    => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready          => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid          => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel        => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data           => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket  => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket    => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			sink2_ready          => rsp_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid          => rsp_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel        => rsp_xbar_demux_002_src0_channel,       --          .channel
			sink2_data           => rsp_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket  => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket    => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink3_ready          => rsp_xbar_demux_003_src0_ready,         --     sink3.ready
			sink3_valid          => rsp_xbar_demux_003_src0_valid,         --          .valid
			sink3_channel        => rsp_xbar_demux_003_src0_channel,       --          .channel
			sink3_data           => rsp_xbar_demux_003_src0_data,          --          .data
			sink3_startofpacket  => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			sink3_endofpacket    => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			sink4_ready          => rsp_xbar_demux_004_src0_ready,         --     sink4.ready
			sink4_valid          => rsp_xbar_demux_004_src0_valid,         --          .valid
			sink4_channel        => rsp_xbar_demux_004_src0_channel,       --          .channel
			sink4_data           => rsp_xbar_demux_004_src0_data,          --          .data
			sink4_startofpacket  => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			sink4_endofpacket    => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			sink5_ready          => rsp_xbar_demux_005_src0_ready,         --     sink5.ready
			sink5_valid          => rsp_xbar_demux_005_src0_valid,         --          .valid
			sink5_channel        => rsp_xbar_demux_005_src0_channel,       --          .channel
			sink5_data           => rsp_xbar_demux_005_src0_data,          --          .data
			sink5_startofpacket  => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			sink5_endofpacket    => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			sink6_ready          => rsp_xbar_demux_006_src0_ready,         --     sink6.ready
			sink6_valid          => rsp_xbar_demux_006_src0_valid,         --          .valid
			sink6_channel        => rsp_xbar_demux_006_src0_channel,       --          .channel
			sink6_data           => rsp_xbar_demux_006_src0_data,          --          .data
			sink6_startofpacket  => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			sink6_endofpacket    => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			sink7_ready          => rsp_xbar_demux_007_src0_ready,         --     sink7.ready
			sink7_valid          => rsp_xbar_demux_007_src0_valid,         --          .valid
			sink7_channel        => rsp_xbar_demux_007_src0_channel,       --          .channel
			sink7_data           => rsp_xbar_demux_007_src0_data,          --          .data
			sink7_startofpacket  => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			sink7_endofpacket    => rsp_xbar_demux_007_src0_endofpacket,   --          .endofpacket
			sink8_ready          => rsp_xbar_demux_008_src0_ready,         --     sink8.ready
			sink8_valid          => rsp_xbar_demux_008_src0_valid,         --          .valid
			sink8_channel        => rsp_xbar_demux_008_src0_channel,       --          .channel
			sink8_data           => rsp_xbar_demux_008_src0_data,          --          .data
			sink8_startofpacket  => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			sink8_endofpacket    => rsp_xbar_demux_008_src0_endofpacket,   --          .endofpacket
			sink9_ready          => rsp_xbar_demux_009_src0_ready,         --     sink9.ready
			sink9_valid          => rsp_xbar_demux_009_src0_valid,         --          .valid
			sink9_channel        => rsp_xbar_demux_009_src0_channel,       --          .channel
			sink9_data           => rsp_xbar_demux_009_src0_data,          --          .data
			sink9_startofpacket  => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			sink9_endofpacket    => rsp_xbar_demux_009_src0_endofpacket,   --          .endofpacket
			sink10_ready         => rsp_xbar_demux_010_src0_ready,         --    sink10.ready
			sink10_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			sink10_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			sink10_data          => rsp_xbar_demux_010_src0_data,          --          .data
			sink10_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			sink10_endofpacket   => rsp_xbar_demux_010_src0_endofpacket,   --          .endofpacket
			sink11_ready         => rsp_xbar_demux_011_src0_ready,         --    sink11.ready
			sink11_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			sink11_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			sink11_data          => rsp_xbar_demux_011_src0_data,          --          .data
			sink11_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			sink11_endofpacket   => rsp_xbar_demux_011_src0_endofpacket,   --          .endofpacket
			sink12_ready         => rsp_xbar_demux_012_src0_ready,         --    sink12.ready
			sink12_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			sink12_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			sink12_data          => rsp_xbar_demux_012_src0_data,          --          .data
			sink12_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			sink12_endofpacket   => rsp_xbar_demux_012_src0_endofpacket,   --          .endofpacket
			sink13_ready         => rsp_xbar_demux_013_src0_ready,         --    sink13.ready
			sink13_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			sink13_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			sink13_data          => rsp_xbar_demux_013_src0_data,          --          .data
			sink13_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			sink13_endofpacket   => rsp_xbar_demux_013_src0_endofpacket,   --          .endofpacket
			sink14_ready         => rsp_xbar_demux_014_src0_ready,         --    sink14.ready
			sink14_valid         => rsp_xbar_demux_014_src0_valid,         --          .valid
			sink14_channel       => rsp_xbar_demux_014_src0_channel,       --          .channel
			sink14_data          => rsp_xbar_demux_014_src0_data,          --          .data
			sink14_startofpacket => rsp_xbar_demux_014_src0_startofpacket, --          .startofpacket
			sink14_endofpacket   => rsp_xbar_demux_014_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_001 : component nios2_ht18_lemonde_streit_rsp_xbar_mux_001
		port map (
			clk                 => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data            => rsp_xbar_mux_001_src_data,             --          .data
			src_channel         => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_003_src1_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_003_src1_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_003_src1_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_003_src1_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_003_src1_endofpacket,   --          .endofpacket
			sink2_ready         => rsp_xbar_demux_013_src1_ready,         --     sink2.ready
			sink2_valid         => rsp_xbar_demux_013_src1_valid,         --          .valid
			sink2_channel       => rsp_xbar_demux_013_src1_channel,       --          .channel
			sink2_data          => rsp_xbar_demux_013_src1_data,          --          .data
			sink2_startofpacket => rsp_xbar_demux_013_src1_startofpacket, --          .startofpacket
			sink2_endofpacket   => rsp_xbar_demux_013_src1_endofpacket,   --          .endofpacket
			sink3_ready         => rsp_xbar_demux_014_src1_ready,         --     sink3.ready
			sink3_valid         => rsp_xbar_demux_014_src1_valid,         --          .valid
			sink3_channel       => rsp_xbar_demux_014_src1_channel,       --          .channel
			sink3_data          => rsp_xbar_demux_014_src1_data,          --          .data
			sink3_startofpacket => rsp_xbar_demux_014_src1_startofpacket, --          .startofpacket
			sink3_endofpacket   => rsp_xbar_demux_014_src1_endofpacket    --          .endofpacket
		);

	width_adapter : component nios2_ht18_lemonde_streit_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 60,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 69,
			IN_PKT_BYTE_CNT_L             => 67,
			IN_PKT_TRANS_COMPRESSED_READ  => 61,
			IN_PKT_BURSTWRAP_H            => 72,
			IN_PKT_BURSTWRAP_L            => 70,
			IN_PKT_BURST_SIZE_H           => 75,
			IN_PKT_BURST_SIZE_L           => 73,
			IN_PKT_RESPONSE_STATUS_H      => 99,
			IN_PKT_RESPONSE_STATUS_L      => 98,
			IN_PKT_TRANS_EXCLUSIVE        => 66,
			IN_PKT_BURST_TYPE_H           => 77,
			IN_PKT_BURST_TYPE_L           => 76,
			IN_ST_DATA_W                  => 100,
			OUT_PKT_ADDR_H                => 42,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 51,
			OUT_PKT_BYTE_CNT_L            => 49,
			OUT_PKT_TRANS_COMPRESSED_READ => 43,
			OUT_PKT_BURST_SIZE_H          => 57,
			OUT_PKT_BURST_SIZE_L          => 55,
			OUT_PKT_RESPONSE_STATUS_H     => 81,
			OUT_PKT_RESPONSE_STATUS_L     => 80,
			OUT_PKT_TRANS_EXCLUSIVE       => 48,
			OUT_PKT_BURST_TYPE_H          => 59,
			OUT_PKT_BURST_TYPE_L          => 58,
			OUT_ST_DATA_W                 => 82,
			ST_CHANNEL_W                  => 15,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => up_clocks_0_sys_clk_clk,            --       clk.clk
			reset                => rst_controller_reset_out_reset,     -- clk_reset.reset
			in_valid             => cmd_xbar_mux_013_src_valid,         --      sink.valid
			in_channel           => cmd_xbar_mux_013_src_channel,       --          .channel
			in_startofpacket     => cmd_xbar_mux_013_src_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_mux_013_src_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_mux_013_src_ready,         --          .ready
			in_data              => cmd_xbar_mux_013_src_data,          --          .data
			out_endofpacket      => width_adapter_src_endofpacket,      --       src.endofpacket
			out_data             => width_adapter_src_data,             --          .data
			out_channel          => width_adapter_src_channel,          --          .channel
			out_valid            => width_adapter_src_valid,            --          .valid
			out_ready            => width_adapter_src_ready,            --          .ready
			out_startofpacket    => width_adapter_src_startofpacket,    --          .startofpacket
			in_command_size_data => "000"                               -- (terminated)
		);

	width_adapter_001 : component nios2_ht18_lemonde_streit_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 42,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 51,
			IN_PKT_BYTE_CNT_L             => 49,
			IN_PKT_TRANS_COMPRESSED_READ  => 43,
			IN_PKT_BURSTWRAP_H            => 54,
			IN_PKT_BURSTWRAP_L            => 52,
			IN_PKT_BURST_SIZE_H           => 57,
			IN_PKT_BURST_SIZE_L           => 55,
			IN_PKT_RESPONSE_STATUS_H      => 81,
			IN_PKT_RESPONSE_STATUS_L      => 80,
			IN_PKT_TRANS_EXCLUSIVE        => 48,
			IN_PKT_BURST_TYPE_H           => 59,
			IN_PKT_BURST_TYPE_L           => 58,
			IN_ST_DATA_W                  => 82,
			OUT_PKT_ADDR_H                => 60,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 69,
			OUT_PKT_BYTE_CNT_L            => 67,
			OUT_PKT_TRANS_COMPRESSED_READ => 61,
			OUT_PKT_BURST_SIZE_H          => 75,
			OUT_PKT_BURST_SIZE_L          => 73,
			OUT_PKT_RESPONSE_STATUS_H     => 99,
			OUT_PKT_RESPONSE_STATUS_L     => 98,
			OUT_PKT_TRANS_EXCLUSIVE       => 66,
			OUT_PKT_BURST_TYPE_H          => 77,
			OUT_PKT_BURST_TYPE_L          => 76,
			OUT_ST_DATA_W                 => 100,
			ST_CHANNEL_W                  => 15,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => up_clocks_0_sys_clk_clk,             --       clk.clk
			reset                => rst_controller_reset_out_reset,      -- clk_reset.reset
			in_valid             => id_router_013_src_valid,             --      sink.valid
			in_channel           => id_router_013_src_channel,           --          .channel
			in_startofpacket     => id_router_013_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_013_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_013_src_ready,             --          .ready
			in_data              => id_router_013_src_data,              --          .data
			out_endofpacket      => width_adapter_001_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_001_src_data,          --          .data
			out_channel          => width_adapter_001_src_channel,       --          .channel
			out_valid            => width_adapter_001_src_valid,         --          .valid
			out_ready            => width_adapter_001_src_ready,         --          .ready
			out_startofpacket    => width_adapter_001_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_002 : component nios2_ht18_lemonde_streit_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 60,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 69,
			IN_PKT_BYTE_CNT_L             => 67,
			IN_PKT_TRANS_COMPRESSED_READ  => 61,
			IN_PKT_BURSTWRAP_H            => 72,
			IN_PKT_BURSTWRAP_L            => 70,
			IN_PKT_BURST_SIZE_H           => 75,
			IN_PKT_BURST_SIZE_L           => 73,
			IN_PKT_RESPONSE_STATUS_H      => 99,
			IN_PKT_RESPONSE_STATUS_L      => 98,
			IN_PKT_TRANS_EXCLUSIVE        => 66,
			IN_PKT_BURST_TYPE_H           => 77,
			IN_PKT_BURST_TYPE_L           => 76,
			IN_ST_DATA_W                  => 100,
			OUT_PKT_ADDR_H                => 42,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 51,
			OUT_PKT_BYTE_CNT_L            => 49,
			OUT_PKT_TRANS_COMPRESSED_READ => 43,
			OUT_PKT_BURST_SIZE_H          => 57,
			OUT_PKT_BURST_SIZE_L          => 55,
			OUT_PKT_RESPONSE_STATUS_H     => 81,
			OUT_PKT_RESPONSE_STATUS_L     => 80,
			OUT_PKT_TRANS_EXCLUSIVE       => 48,
			OUT_PKT_BURST_TYPE_H          => 59,
			OUT_PKT_BURST_TYPE_L          => 58,
			OUT_ST_DATA_W                 => 82,
			ST_CHANNEL_W                  => 15,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => up_clocks_0_sys_clk_clk,             --       clk.clk
			reset                => rst_controller_reset_out_reset,      -- clk_reset.reset
			in_valid             => cmd_xbar_mux_014_src_valid,          --      sink.valid
			in_channel           => cmd_xbar_mux_014_src_channel,        --          .channel
			in_startofpacket     => cmd_xbar_mux_014_src_startofpacket,  --          .startofpacket
			in_endofpacket       => cmd_xbar_mux_014_src_endofpacket,    --          .endofpacket
			in_ready             => cmd_xbar_mux_014_src_ready,          --          .ready
			in_data              => cmd_xbar_mux_014_src_data,           --          .data
			out_endofpacket      => width_adapter_002_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_002_src_data,          --          .data
			out_channel          => width_adapter_002_src_channel,       --          .channel
			out_valid            => width_adapter_002_src_valid,         --          .valid
			out_ready            => width_adapter_002_src_ready,         --          .ready
			out_startofpacket    => width_adapter_002_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_003 : component nios2_ht18_lemonde_streit_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 42,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 51,
			IN_PKT_BYTE_CNT_L             => 49,
			IN_PKT_TRANS_COMPRESSED_READ  => 43,
			IN_PKT_BURSTWRAP_H            => 54,
			IN_PKT_BURSTWRAP_L            => 52,
			IN_PKT_BURST_SIZE_H           => 57,
			IN_PKT_BURST_SIZE_L           => 55,
			IN_PKT_RESPONSE_STATUS_H      => 81,
			IN_PKT_RESPONSE_STATUS_L      => 80,
			IN_PKT_TRANS_EXCLUSIVE        => 48,
			IN_PKT_BURST_TYPE_H           => 59,
			IN_PKT_BURST_TYPE_L           => 58,
			IN_ST_DATA_W                  => 82,
			OUT_PKT_ADDR_H                => 60,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 69,
			OUT_PKT_BYTE_CNT_L            => 67,
			OUT_PKT_TRANS_COMPRESSED_READ => 61,
			OUT_PKT_BURST_SIZE_H          => 75,
			OUT_PKT_BURST_SIZE_L          => 73,
			OUT_PKT_RESPONSE_STATUS_H     => 99,
			OUT_PKT_RESPONSE_STATUS_L     => 98,
			OUT_PKT_TRANS_EXCLUSIVE       => 66,
			OUT_PKT_BURST_TYPE_H          => 77,
			OUT_PKT_BURST_TYPE_L          => 76,
			OUT_ST_DATA_W                 => 100,
			ST_CHANNEL_W                  => 15,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => up_clocks_0_sys_clk_clk,             --       clk.clk
			reset                => rst_controller_reset_out_reset,      -- clk_reset.reset
			in_valid             => id_router_014_src_valid,             --      sink.valid
			in_channel           => id_router_014_src_channel,           --          .channel
			in_startofpacket     => id_router_014_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_014_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_014_src_ready,             --          .ready
			in_data              => id_router_014_src_data,              --          .data
			out_endofpacket      => width_adapter_003_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_003_src_data,          --          .data
			out_channel          => width_adapter_003_src_channel,       --          .channel
			out_valid            => width_adapter_003_src_valid,         --          .valid
			out_ready            => width_adapter_003_src_ready,         --          .ready
			out_startofpacket    => width_adapter_003_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	irq_mapper : component nios2_ht18_lemonde_streit_irq_mapper
		port map (
			clk           => up_clocks_0_sys_clk_clk,             --       clk.clk
			reset         => rst_controller_reset_out_reset,      -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,            -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,            -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,            -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,            -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,            -- receiver4.irq
			sender_irq    => nios2_ht18_lemonde_streit_d_irq_irq  --    sender.irq
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv <= not jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;

	jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv <= not jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;

	timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv <= not timer_0_s1_translator_avalon_anti_slave_0_write;

	timer_1_s1_translator_avalon_anti_slave_0_write_ports_inv <= not timer_1_s1_translator_avalon_anti_slave_0_write;

	de2_pio_toggles18_s1_translator_avalon_anti_slave_0_write_ports_inv <= not de2_pio_toggles18_s1_translator_avalon_anti_slave_0_write;

	de2_pio_keys4_s1_translator_avalon_anti_slave_0_write_ports_inv <= not de2_pio_keys4_s1_translator_avalon_anti_slave_0_write;

	de2_pio_redled18_s1_translator_avalon_anti_slave_0_write_ports_inv <= not de2_pio_redled18_s1_translator_avalon_anti_slave_0_write;

	de2_pio_greenled9_s1_translator_avalon_anti_slave_0_write_ports_inv <= not de2_pio_greenled9_s1_translator_avalon_anti_slave_0_write;

	de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_write_ports_inv <= not de2_pio_hex_high28_s1_translator_avalon_anti_slave_0_write;

	de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_write_ports_inv <= not de2_pio_hex_low28_s1_translator_avalon_anti_slave_0_write;

	sdram_s1_translator_avalon_anti_slave_0_write_ports_inv <= not sdram_s1_translator_avalon_anti_slave_0_write;

	sdram_s1_translator_avalon_anti_slave_0_read_ports_inv <= not sdram_s1_translator_avalon_anti_slave_0_read;

	sdram_s1_translator_avalon_anti_slave_0_byteenable_ports_inv <= not sdram_s1_translator_avalon_anti_slave_0_byteenable;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of nios2_ht18_lemonde_streit
